//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "new.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "coke"
//: require "74xxGateLevel"
//: require "tty"
//: require "m68xx"
//: require "timer"
//: require "74xx"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w58;    //: /sn:0 {0}(794,982)(776,982)(776,936)(759,936){1}
reg w50;    //: /sn:0 {0}(480,-318)(460,-318)(460,-116)(424,-116){1}
reg w72;    //: /sn:0 {0}(318,-341)(318,-326)(275,-326){1}
reg w22;    //: /sn:0 {0}(702,208)(724,208)(724,208)(751,208){1}
reg w20;    //: /sn:0 {0}(332,-95)(332,-184){1}
reg w18;    //: /sn:0 {0}(556,-323)(619,-323){1}
supply0 w19;    //: /sn:0 {0}(339,-261)(339,-234){1}
supply0 w23;    //: /sn:0 {0}(292,-302)(292,-316)(275,-316){1}
reg w54;    //: /sn:0 {0}(870,977)(969,977)(969,960){1}
reg w24;    //: /sn:0 {0}(702,258)(724,258)(724,258)(751,258){1}
reg [7:0] w31;    //: /sn:0 {0}(#:209,-599)(209,-577)(220,-577)(220,-562){1}
reg w53;    //: /sn:0 {0}(660,394)(788,394){1}
//: {2}(792,394)(979,394)(979,448)(962,448){3}
//: {4}(790,396)(790,449)(775,449){5}
supply0 w46;    //: /sn:0 {0}(979,476)(979,458)(962,458){1}
reg w8;    //: /sn:0 {0}(132,-321)(211,-321)(211,-321)(199,-321){1}
reg w52;    //: /sn:0 {0}(661,454)(677,454){1}
//: {2}(681,454)(699,454){3}
//: {4}(679,452)(679,421)(871,421)(871,453)(886,453){5}
supply1 w17;    //: /sn:0 {0}(363,-159)(346,-159)(346,-184){1}
supply0 w27;    //: /sn:0 {0}(260,-548)(276,-548)(276,-511)(293,-511){1}
supply0 w47;    //: /sn:0 {0}(887,1023)(887,987)(870,987){1}
supply1 w76;    //: /sn:0 {0}(352,997)(379,997)(379,978)(430,978){1}
supply0 w26;    //: /sn:0 {0}(556,-313)(571,-313)(571,-296){1}
supply0 w51;    //: /sn:0 {0}(792,473)(792,459)(775,459){1}
wire [15:0] w16;    //: /sn:0 {0}(#:517,-307)(517,-278){1}
//: {2}(#:519,-276)(743,-276)(743,-311){3}
//: {4}(517,-274)(517,-223){5}
//: {6}(517,-222)(517,-199){7}
//: {8}(517,-198)(517,-179){9}
//: {10}(517,-178)(517,-139){11}
//: {12}(517,-138)(517,-55){13}
//: {14}(517,-54)(517,-30){15}
//: {16}(517,-29)(517,14){17}
//: {18}(517,15)(517,40){19}
//: {20}(517,41)(517,58){21}
wire [7:0] w13;    //: /sn:0 {0}(#:736,444)(736,382){1}
//: {2}(738,380)(1442,380)(1442,750)(1405,750){3}
//: {4}(736,378)(736,365){5}
//: {6}(736,361)(736,345)(#:772,345)(#:772,332){7}
//: {8}(#:734,363)(667,363)(667,335){9}
wire [7:0] w6;    //: /sn:0 {0}(#:832,891)(832,937){1}
//: {2}(#:834,939)(879,939)(879,925){3}
//: {4}(832,941)(832,948)(831,948)(831,972){5}
wire [7:0] w65;    //: /sn:0 {0}(#:1495,851)(1506,851)(1506,851)(1549,851)(1549,715)(1571,715){1}
//: {2}(1573,713)(1573,-312){3}
//: {4}(1573,-316)(1573,-474)(842,-474)(#:842,-399){5}
//: {6}(#:1571,-314)(1472,-314)(1472,-347){7}
//: {8}(1573,717)(1573,718)(1640,718)(#:1640,656){9}
wire w7;    //: /sn:0 {0}(402,301)(407,301){1}
//: {2}(411,301)(439,301){3}
//: {4}(443,301)(453,301)(453,87)(712,87){5}
//: {6}(716,87)(751,87){7}
//: {8}(714,85)(714,78)(714,78)(714,72){9}
//: {10}(441,299)(441,275){11}
//: {12}(409,303)(409,968)(430,968){13}
wire w34;    //: /sn:0 {0}(356,858)(34,858)(34,443){1}
//: {2}(36,441)(119,441){3}
//: {4}(123,441)(202,441)(202,306)(381,306){5}
//: {6}(121,443)(121,576)(379,576){7}
//: {8}(32,441)(-24,441)(-24,441)(-66,441){9}
//: {10}(-68,439)(-68,436)(-68,436)(-68,426){11}
//: {12}(-70,441)(-80,441)(-80,441)(-75,441){13}
wire w81;    //: /sn:0 {0}(-83,-261)(-83,-35)(-48,-35)(-48,48){1}
//: {2}(-46,50)(-54,50)(-54,50)(-12,50){3}
//: {4}(-50,50)(-66,50)(-66,50)(-75,50){5}
wire [7:0] w59;    //: /sn:0 {0}(#:832,-370)(832,-347)(832,-347)(832,-322){1}
//: {2}(834,-320)(946,-320)(946,-346){3}
//: {4}(832,-318)(#:832,-104){5}
wire w25;    //: /sn:0 {0}(737,1225)(737,1199)(737,1199)(737,1054){1}
//: {2}(739,1052)(815,1052)(815,1036){3}
//: {4}(737,1050)(737,1018)(516,1018){5}
wire [7:0] w62;    //: /sn:0 {0}(#:1225,788)(1192,788){1}
//: {2}(1190,786)(#:1190,780)(1190,780)(1190,718){3}
//: {4}(1188,788)(1154,788)(1154,-198)(970,-198){5}
//: {6}(968,-200)(968,-275){7}
//: {8}(966,-198)(521,-198){9}
wire w39;    //: /sn:0 {0}(-75,228)(-68,228){1}
//: {2}(-64,228)(189,228)(189,286)(381,286){3}
//: {4}(-66,226)(-66,210){5}
wire [7:0] w4;    //: /sn:0 {0}(#:746,598)(746,632){1}
//: {2}(748,634)(1375,634)(#:1375,502){3}
//: {4}(746,636)(746,663){5}
//: {6}(#:744,665)(686,665)(686,640){7}
//: {8}(746,667)(746,691)(786,691)(786,704){9}
wire w56;    //: /sn:0 {0}(-68,526)(-68,550)(-68,550)(-68,533){1}
//: {2}(-66,535)(50,535){3}
//: {4}(54,535)(158,535){5}
//: {6}(162,535)(219,535)(219,321)(381,321){7}
//: {8}(160,537)(160,591)(379,591){9}
//: {10}(52,537)(52,873)(356,873){11}
//: {12}(-70,535)(-75,535){13}
wire [7:0] w0;    //: /sn:0 {0}(#:99,-635)(139,-635)(139,-671)(221,-671){1}
//: {2}(225,-671)(#:252,-671)(252,-562){3}
//: {4}(223,-673)(223,-717){5}
wire [7:0] w3;    //: /sn:0 {0}(#:831,993)(831,1040){1}
//: {2}(833,1042)(922,1042)(922,1019){3}
//: {4}(#:831,1044)(831,1242)(787,1242){5}
wire w36;    //: /sn:0 {0}(381,296)(190,296)(190,361)(25,361){1}
//: {2}(21,361)(0,361){3}
//: {4}(-4,361)(-63,361){5}
//: {6}(-65,359)(-65,343){7}
//: {8}(-67,361)(-75,361){9}
//: {10}(-2,363)(-2,1021)(424,1021)(424,1020)(495,1020){11}
//: {12}(23,363)(23,848)(356,848){13}
wire [7:0] w60;    //: /sn:0 {0}(#:943,569)(943,558){1}
//: {2}(#:945,556)(988,556)(988,545){3}
//: {4}(943,554)(943,516)(1284,516)(1284,-222)(1063,-222){5}
//: {6}(1061,-224)(1061,-276){7}
//: {8}(1059,-222)(521,-222){9}
wire [3:0] w29;    //: /sn:0 {0}(#:-266,25)(-315,25)(-315,-49)(-130,-49){1}
//: {2}(-126,-49)(146,-49)(146,41)(427,41){3}
//: {4}(431,41)(443,41){5}
//: {6}(447,41)(512,41){7}
//: {8}(445,39)(#:445,40)(445,40)(445,-24){9}
//: {10}(429,43)(429,797)(666,797){11}
//: {12}(670,797)(#:707,797){13}
//: {14}(668,795)(668,792)(668,792)(668,760){15}
//: {16}(#:-128,-51)(-128,-107){17}
wire w30;    //: /sn:0 {0}(-75,312)(-69,312){1}
//: {2}(-65,312)(16,312){3}
//: {4}(20,312)(55,312)(55,312)(82,312){5}
//: {6}(86,312)(186,312)(186,291)(381,291){7}
//: {8}(84,314)(84,566)(379,566){9}
//: {10}(18,314)(18,487)(132,487)(132,843)(356,843){11}
//: {12}(-67,310)(-67,292){13}
wire w71;    //: /sn:0 {0}(377,855)(390,855){1}
//: {2}(394,855)(492,855){3}
//: {4}(496,855)(591,855)(591,149)(644,149){5}
//: {6}(648,149)(751,149){7}
//: {8}(646,147)(646,137)(646,137)(646,71){9}
//: {10}(494,853)(494,841){11}
//: {12}(392,857)(392,973)(430,973){13}
wire [7:0] w37;    //: /sn:0 {0}(#:923,464)(923,491){1}
//: {2}(#:925,493)(1021,493)(1021,477){3}
//: {4}(923,495)(923,569){5}
wire [2:0] w12;    //: /sn:0 {0}(#:908,34)(936,34){1}
//: {2}(940,34)(#:1014,34){3}
//: {4}(938,32)(#:938,38)(938,38)(938,12){5}
wire w73;    //: /sn:0 {0}(809,-383)(776,-383)(776,-333)(968,-333)(968,-35){1}
//: {2}(970,-33)(987,-33){3}
//: {4}(991,-33)(1027,-33)(1027,11){5}
//: {6}(989,-35)(989,-45)(989,-45)(989,-55){7}
//: {8}(966,-33)(961,-33)(961,290)(1091,290)(1091,742){9}
//: {10}(1093,744)(1241,744){11}
//: {12}(1245,744)(1369,744)(1369,772)(1440,772)(1440,834)(1487,834)(1487,846){13}
//: {14}(1243,746)(1243,763){15}
//: {16}(1089,744)(1061,744){17}
//: {18}(1057,744)(1025,744){19}
//: {20}(1021,744)(949,744){21}
//: {22}(1023,746)(1023,754)(1023,754)(1023,730){23}
//: {24}(1059,746)(1059,790)(1080,790){25}
wire [2:0] w10;    //: /sn:0 {0}(#:1043,44)(1071,44)(1071,-138)(617,-138){1}
//: {2}(615,-140)(#:615,-149)(615,-149)(615,-251){3}
//: {4}(613,-138)(521,-138){5}
wire w70;    //: /sn:0 {0}(150,-532)(184,-532)(184,-548)(212,-548){1}
wire [15:0] w21;    //: /sn:0 {0}(517,-328)(517,-347)(#:426,-347)(426,-211)(373,-211){1}
//: {2}(371,-213)(#:371,-223)(371,-223)(371,-298){3}
//: {4}(369,-211)(#:356,-211){5}
wire [2:0] w1;    //: /sn:0 {0}(#:751,-29)(639,-29){1}
//: {2}(637,-31)(637,-82){3}
//: {4}(635,-29)(521,-29){5}
wire w68;    //: /sn:0 {0}(451,973)(476,973)(476,1015)(495,1015){1}
wire w32;    //: /sn:0 {0}(356,868)(46,868)(46,508){1}
//: {2}(48,506)(168,506){3}
//: {4}(172,506)(213,506)(213,316)(381,316){5}
//: {6}(170,508)(170,586)(379,586){7}
//: {8}(44,506)(-12,506)(-12,506)(-67,506){9}
//: {10}(-69,504)(-69,498)(-69,498)(-69,493){11}
//: {12}(-71,506)(-73,506)(-73,506)(-75,506){13}
wire w44;    //: /sn:0 {0}(-10,117)(-56,117)(-56,117)(-55,117){1}
//: {2}(-57,115)(-57,-22)(-93,-22)(-93,-261){3}
//: {4}(-59,117)(-63,117)(-63,117)(-75,117){5}
wire [7:0] w75;    //: /sn:0 {0}(#:673,1251)(-584,1251)(-584,-645)(70,-645){1}
wire w35;    //: /sn:0 {0}(356,853)(28,853)(28,409){1}
//: {2}(30,407)(107,407){3}
//: {4}(111,407)(197,407)(197,301)(381,301){5}
//: {6}(109,409)(109,571)(379,571){7}
//: {8}(26,407)(-64,407){9}
//: {10}(-66,405)(-66,402)(-66,402)(-66,392){11}
//: {12}(-68,407)(-75,407){13}
wire w33;    //: /sn:0 {0}(356,863)(40,863)(40,474){1}
//: {2}(42,472)(83,472)(83,472)(129,472){3}
//: {4}(133,472)(208,472)(208,311)(381,311){5}
//: {6}(131,474)(131,581)(379,581){7}
//: {8}(38,472)(-18,472)(-18,472)(-67,472){9}
//: {10}(-69,470)(-69,466)(-69,466)(-69,459){11}
//: {12}(-71,472)(-77,472)(-77,472)(-75,472){13}
wire [7:0] w28;    //: /sn:0 {0}(#:236,-331)(236,-392){1}
//: {2}(#:238,-394)(331,-394)(331,-402){3}
//: {4}(236,-396)(#:236,-533){5}
wire w49;    //: /sn:0 {0}(949,799)(959,799)(959,799)(964,799){1}
wire w45;    //: /sn:0 {0}(-78,-261)(-78,-42)(-43,-42)(-43,15){1}
//: {2}(-41,17)(-54,17)(-54,17)(-14,17){3}
//: {4}(-45,17)(-63,17)(-63,17)(-75,17){5}
wire [7:0] w14;    //: /sn:0 {0}(#:923,443)(923,365){1}
//: {2}(#:925,363)(970,363)(970,336){3}
//: {4}(923,361)(923,341)(886,341)(#:886,332){5}
wire w69;    //: /sn:0 {0}(1026,874)(1026,862){1}
//: {2}(1028,860)(1057,860){3}
//: {4}(1061,860)(1250,860)(1250,835){5}
//: {6}(1252,833)(1397,833)(1397,755){7}
//: {8}(1250,831)(1250,813){9}
//: {10}(1059,858)(1059,795)(1080,795){11}
//: {12}(1026,858)(1026,857)(949,857){13}
wire [7:0] w48;    //: /sn:0 {0}(#:1260,786)(1305,786){1}
//: {2}(1309,786)(1318,786){3}
//: {4}(1322,786)(1414,786)(1414,851)(1479,851){5}
//: {6}(1320,788)(1320,804)(1320,804)(1320,850){7}
//: {8}(1307,784)(1307,750)(#:1389,750){9}
wire w78;    //: /sn:0 {0}(1101,793)(1213,793)(1213,837)(1236,837)(1236,813){1}
wire [2:0] w11;    //: /sn:0 {0}(#:1043,24)(1114,24)(1114,-178)(897,-178){1}
//: {2}(895,-180)(#:895,-257){3}
//: {4}(893,-178)(521,-178){5}
wire w41;    //: /sn:0 {0}(-75,157)(-66,157){1}
//: {2}(-62,157)(59,157){3}
//: {4}(63,157)(196,157)(196,276)(381,276){5}
//: {6}(61,159)(61,561)(379,561){7}
//: {8}(-64,155)(-64,144){9}
wire [2:0] w2;    //: /sn:0 {0}(#:751,15)(732,15){1}
//: {2}(730,13)(730,-80){3}
//: {4}(728,15)(521,15){5}
wire [7:0] w85;    //: /sn:0 {0}(#:673,1296)(-483,1296)(-483,-475)(822,-475)(#:822,-399){1}
wire [7:0] w15;    //: /sn:0 {0}(#:236,-310)(236,-269){1}
//: {2}(234,-267)(55,-267)(55,-625)(70,-625){3}
//: {4}(236,-265)(236,-247){5}
//: {6}(#:234,-245)(22,-245)(22,-268){7}
//: {8}(236,-243)(236,-221)(237,-221)(237,-211){9}
//: {10}(239,-209)(274,-209){11}
//: {12}(278,-209)(321,-209){13}
//: {14}(276,-211)(276,-253){15}
//: {16}(237,-207)(237,518)(756,518)(756,551){17}
//: {18}(#:754,553)(671,553)(671,543){19}
//: {20}(756,555)(756,569){21}
wire w55;    //: /sn:0 {0}(569,1038)(569,1054)(609,1054){1}
//: {2}(613,1054)(709,1054)(709,1225){3}
//: {4}(611,1052)(611,587){5}
//: {6}(613,585)(632,585){7}
//: {8}(636,585)(723,585){9}
//: {10}(634,587)(634,646)(907,646)(907,585)(910,585){11}
//: {12}(609,585)(483,585)(483,-54)(512,-54){13}
wire w38;    //: /sn:0 {0}(-75,271)(-74,271)(-74,271)(-70,271){1}
//: {2}(-66,271)(12,271)(12,838)(356,838){3}
//: {4}(-68,269)(-68,259)(-68,259)(-68,250){5}
wire [7:0] w5;    //: /sn:0 {0}(#:933,598)(933,670){1}
//: {2}(#:935,672)(1004,672)(1004,659){3}
//: {4}(933,674)(933,691)(894,691)(#:894,704){5}
wire w43;    //: /sn:0 {0}(-88,-261)(-88,-29)(-52,-29)(-52,79){1}
//: {2}(-50,81)(-54,81)(-54,81)(-10,81){3}
//: {4}(-54,81)(-75,81){5}
wire w64;    //: /sn:0 {0}(400,578)(451,578){1}
//: {2}(455,578)(549,578)(549,120)(675,120){3}
//: {4}(679,120)(751,120){5}
//: {6}(677,118)(677,93)(677,93)(677,72){7}
//: {8}(453,576)(453,571)(453,571)(453,559){9}
wire [7:0] w9;    //: /sn:0 {0}(#:736,465)(736,500){1}
//: {2}(#:734,502)(641,502)(641,487){3}
//: {4}(736,504)(736,569){5}
wire w77;    //: /sn:0 {0}(-86,-282)(-86,-597)(86,-597)(86,-612){1}
wire w57;    //: /sn:0 {0}(356,878)(58,878)(58,566){1}
//: {2}(60,564)(150,564){3}
//: {4}(154,564)(224,564)(224,326)(381,326){5}
//: {6}(152,566)(152,596)(379,596){7}
//: {8}(56,564)(-65,564){9}
//: {10}(-67,562)(-67,555){11}
//: {12}(-69,564)(-75,564){13}
wire w40;    //: /sn:0 {0}(381,281)(192,281)(192,191)(8,191){1}
//: {2}(4,191)(-35,191)(-35,191)(-60,191){3}
//: {4}(-62,189)(-62,183)(-62,183)(-62,173){5}
//: {6}(-64,191)(-77,191)(-77,191)(-75,191){7}
//: {8}(6,193)(6,833)(356,833){9}
//: enddecls

  //: LED g164 (w12) @(938,5) /sn:0 /w:[ 5 ] /type:1
  //: GROUND g8 (w26) @(571,-290) /sn:0 /w:[ 1 ]
  //: VDD g4 (w17) @(363,-148) /sn:0 /R:3 /w:[ 0 ]
  //: DIP g116 (w31) @(209,-609) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: LED g197 (w71) @(646,64) /sn:0 /w:[ 9 ] /type:0
  //: joint g157 (w25) @(737, 1052) /w:[ 2 4 -1 1 ]
  assign w10 = w16[11:9]; //: TAP g17 @(515,-138) /sn:0 /R:2 /w:[ 5 12 11 ] /ss:1
  //: LED g137 (w45) @(-7,17) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: LED g74 (w48) @(1320,857) /sn:0 /R:2 /w:[ 7 ] /type:1
  //: joint g198 (w71) @(646, 149) /w:[ 6 8 5 -1 ]
  //: joint g30 (w57) @(58, 564) /w:[ 2 -1 8 1 ]
  //: joint g92 (w6) @(832, 939) /w:[ 2 1 -1 4 ]
  //: joint g77 (w48) @(1320, 786) /w:[ 4 -1 3 6 ]
  //: joint g130 (w62) @(968, -198) /w:[ 5 6 8 -1 ]
  _GGREG8 #(10, 10, 20) PC (.Q(w15), .D(w28), .EN(w23), .CLR(~w72), .CK(w8));   //: @(236,-321) /w:[ 0 0 1 1 1 ]
  _GGRAM8x16 #(10, 60, 70, 10, 10, 10) g1 (.A(w15), .D(w21), .WE(~w19), .OE(~w17), .CS(~w20));   //: @(339,-210) /sn:0 /w:[ 13 5 1 1 1 ]
  //: joint g214 (w48) @(1307, 786) /w:[ 2 8 1 -1 ]
  //: joint g111 (w65) @(1573, -314) /w:[ -1 4 6 3 ]
  //: LED g179 (w30) @(-67,285) /sn:0 /w:[ 13 ] /type:0
  //: joint g144 (w4) @(746, 665) /w:[ -1 5 6 8 ]
  assign w60 = w16[11:4]; //: TAP g51 @(515,-222) /sn:0 /R:2 /w:[ 9 6 5 ] /ss:1
  //: joint g70 (w33) @(-69, 472) /w:[ 9 10 12 -1 ]
  //: joint g161 (w64) @(453, 578) /w:[ 2 8 1 -1 ]
  //: LED g149 (w62) @(1190,711) /sn:0 /w:[ 3 ] /type:1
  //: joint g25 (w34) @(121, 441) /w:[ 4 -1 3 6 ]
  //: SWITCH g10 (w22) @(685,208) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g65 (w36) @(-2, 361) /w:[ 3 -1 4 10 ]
  //: LED g103 (w16) @(743,-318) /sn:0 /w:[ 3 ] /type:1
  //: joint g64 (w71) @(392, 855) /w:[ 2 -1 1 12 ]
  //: joint g72 (w65) @(1573, 715) /w:[ -1 2 1 8 ]
  //: joint g49 (w15) @(237, -209) /w:[ 10 9 -1 16 ]
  //: SWITCH g6 (w72) @(318,-354) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: joint g142 (w29) @(668, 797) /w:[ 12 14 11 -1 ]
  //: joint g136 (w29) @(445, 41) /w:[ 6 8 5 -1 ]
  //: SWITCH g58 (w58) @(742,936) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: GROUND g56 (w47) @(887,1029) /sn:0 /w:[ 0 ]
  //: joint g35 (w35) @(28, 407) /w:[ 2 -1 8 1 ]
  //: GROUND g7 (w23) @(292,-296) /sn:0 /w:[ 0 ]
  //: joint g124 (w1) @(637, -29) /w:[ 1 2 4 -1 ]
  //: joint g98 (w30) @(-67, 312) /w:[ 2 12 1 -1 ]
  //: joint g200 (w13) @(736, 380) /w:[ 2 4 -1 1 ]
  //: LED g181 (w36) @(-65,336) /sn:0 /w:[ 7 ] /type:0
  //: joint g67 (w57) @(-67, 564) /w:[ 9 10 12 -1 ]
  //: LED g85 (w9) @(641,480) /sn:0 /w:[ 3 ] /type:1
  //: joint g126 (w2) @(730, 15) /w:[ 1 2 4 -1 ]
  _GGOR2 #(6) g208 (.I0(w68), .I1(w36), .Z(w25));   //: @(506,1018) /sn:0 /w:[ 1 11 5 ]
  assign w29 = w16[15:12]; //: TAP g54 @(515,41) /sn:0 /R:2 /w:[ 7 20 19 ] /ss:0
  //: joint g33 (w33) @(40, 472) /w:[ 2 -1 8 1 ]
  //: joint g52 (w41) @(-64, 157) /w:[ 2 8 1 -1 ]
  //: joint g40 (w44) @(-57, 117) /w:[ 1 2 4 -1 ]
  _GGREG8 #(10, 10, 20) RA (.Q(w9), .D(w13), .EN(w51), .CLR(~w53), .CK(w52));   //: @(736,454) /w:[ 0 0 1 5 3 ]
  //: LED g81 (w13) @(667,328) /sn:0 /w:[ 9 ] /type:1
  //: joint g163 (w7) @(441, 301) /w:[ 4 10 3 -1 ]
  //: joint g132 (w11) @(895, -178) /w:[ 1 2 4 -1 ]
  _GGOR2 #(6) g210 (.I0(w73), .I1(w69), .Z(w78));   //: @(1091,793) /sn:0 /w:[ 25 11 0 ]
  assign w1 = w16[11:9]; //: TAP g12 @(515,-29) /sn:0 /R:2 /w:[ 5 16 15 ] /ss:1
  //: LED g108 (w59) @(946,-353) /sn:0 /w:[ 3 ] /type:1
  _GGBUFIF8 #(4, 6) g106 (.Z(w48), .I(w13), .E(w69));   //: @(1399,750) /sn:0 /R:2 /w:[ 9 3 7 ]
  //: LED g131 (w11) @(895,-264) /sn:0 /w:[ 3 ] /type:1
  //: joint g194 (w7) @(714, 87) /w:[ 6 8 5 -1 ]
  //: LED g177 (w38) @(-68,243) /sn:0 /w:[ 5 ] /type:0
  //: joint g96 (w35) @(-66, 407) /w:[ 9 10 12 -1 ]
  _GGREG8 #(10, 10, 20) RB (.Q(w37), .D(w14), .EN(w46), .CLR(~w53), .CK(w52));   //: @(923,453) /w:[ 0 0 1 3 5 ]
  //: VDD g209 (w76) @(352,986) /sn:0 /R:1 /w:[ 0 ]
  //: joint g196 (w64) @(677, 120) /w:[ 4 6 3 -1 ]
  ALU g19 (.RA(w4), .RB(w5), .ALU_op(w29), .ALU_OUTPUT(w6), .LOAD(w73), .MOV(w49), .STR(w69));   //: @(708, 705) /sz:(240, 185) /R:3 /sn:0 /p:[ Ti0>9 Ti1>5 Li0>13 Bo0<0 Ro0<21 Ro1<0 Ro2<13 ]
  _GGADD8 #(68, 70, 62, 64) g114 (.A(w31), .B(w0), .S(w28), .CI(w27), .CO(w70));   //: @(236,-546) /sn:0 /w:[ 1 3 5 0 1 ]
  //: LED g117 (w70) @(143,-532) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: joint g78 (w15) @(236, -245) /w:[ -1 5 6 8 ]
  //: LED g125 (w2) @(730,-87) /sn:0 /w:[ 3 ] /type:1
  //: joint g155 (w39) @(-66, 228) /w:[ 2 4 1 -1 ]
  _GGMUX2x8 #(8, 8) g105 (.I0(w85), .I1(w65), .S(w73), .Z(w59));   //: @(832,-383) /sn:0 /w:[ 1 5 0 0 ] /ss:0 /do:0
  //: joint g63 (w7) @(409, 301) /w:[ 2 -1 1 12 ]
  //: LED g93 (w3) @(922,1012) /sn:0 /w:[ 3 ] /type:1
  //: joint g100 (w73) @(1023, 744) /w:[ 19 -1 20 22 ]
  //: SWITCH g113 (w8) @(115,-321) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g212 (w69) @(1059, 860) /w:[ 4 10 3 -1 ]
  //: joint g211 (w73) @(1059, 744) /w:[ 17 -1 18 24 ]
  //: GROUND g43 (w51) @(792,479) /sn:0 /w:[ 0 ]
  //: joint g38 (w40) @(6, 191) /w:[ 1 -1 2 8 ]
  register_file g0 (.C(w59), .CLR(w24), .CLK(w22), .rc_s(w71), .rb_s(w64), .ra_s(w7), .Add_B(w2), .Add_A(w1), .Add_C(w12), .B(w14), .A(w13));   //: @(752, -103) /sz:(155, 434) /sn:0 /p:[ Ti0>5 Li0>1 Li1>1 Li2>7 Li3>5 Li4>7 Li5>0 Li6>0 Ri0>0 Bo0<5 Bo1<7 ]
  //: LED g101 (w69) @(1026,881) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g48 (w45) @(-43, 17) /w:[ 2 1 4 -1 ]
  _GGREG8 #(10, 10, 20) RZ (.Q(w3), .D(w6), .EN(w47), .CLR(~w54), .CK(w58));   //: @(831,982) /w:[ 0 5 1 0 0 ]
  //: joint g37 (w30) @(18, 312) /w:[ 4 -1 3 10 ]
  //: joint g95 (w34) @(-68, 441) /w:[ 9 10 12 -1 ]
  //: joint g80 (w14) @(923, 363) /w:[ 2 4 -1 1 ]
  //: LED g120 (w15) @(276,-260) /sn:0 /w:[ 15 ] /type:1
  //: joint g122 (w21) @(371, -211) /w:[ 1 2 4 -1 ]
  //: LED g76 (w15) @(22,-275) /sn:0 /w:[ 7 ] /type:1
  //: LED g189 (w56) @(-68,519) /sn:0 /w:[ 0 ] /type:0
  //: LED g170 (w0) @(223,-724) /sn:0 /w:[ 5 ] /type:1
  //: LED g152 (w65) @(1640,649) /sn:0 /w:[ 9 ] /type:1
  assign w62 = w16[8:1]; //: TAP g75 @(515,-198) /sn:0 /R:2 /w:[ 9 8 7 ] /ss:1
  //: GROUND g44 (w46) @(979,482) /sn:0 /w:[ 0 ]
  //: joint g47 (w81) @(-48, 50) /w:[ 2 1 4 -1 ]
  //: LED g182 (w35) @(-66,385) /sn:0 /w:[ 11 ] /type:0
  //: joint g159 (w71) @(494, 855) /w:[ 4 10 3 -1 ]
  assign w11 = w16[5:3]; //: TAP g16 @(515,-178) /sn:0 /R:2 /w:[ 5 10 9 ] /ss:1
  //: GROUND g3 (w19) @(339,-267) /sn:0 /R:2 /w:[ 0 ]
  //: joint g109 (w73) @(968, -33) /w:[ 2 1 8 -1 ]
  //: LED g143 (w4) @(686,633) /sn:0 /w:[ 7 ] /type:1
  //: joint g26 (w35) @(109, 407) /w:[ 4 -1 3 6 ]
  _GGREG16 #(10, 10, 20) IR (.Q(w16), .D(w21), .EN(w26), .CLR(~w18), .CK(w50));   //: @(517,-318) /w:[ 0 0 0 0 0 ]
  //: joint g90 (w15) @(756, 553) /w:[ -1 17 18 20 ]
  //: LED g174 (w40) @(-62,166) /sn:0 /w:[ 5 ] /type:0
  //: LED g158 (w71) @(494,834) /sn:0 /w:[ 11 ] /type:0
  //: joint g128 (w60) @(1061, -222) /w:[ 5 6 8 -1 ]
  //: SWITCH g2 (w20) @(332,-81) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:1
  //: joint g23 (w32) @(170, 506) /w:[ 4 -1 3 6 ]
  //: LED g91 (w6) @(879,918) /sn:0 /w:[ 3 ] /type:1
  //: joint g39 (w43) @(-52, 81) /w:[ 2 1 4 -1 ]
  //: LED g141 (w29) @(668,753) /sn:0 /w:[ 15 ] /type:1
  //: LED g127 (w60) @(1061,-283) /sn:0 /w:[ 7 ] /type:1
  //: joint g24 (w33) @(131, 472) /w:[ 4 -1 3 6 ]
  //: joint g86 (w9) @(736, 502) /w:[ -1 1 2 4 ]
  //: joint g104 (w16) @(517, -276) /w:[ 2 1 -1 4 ]
  //: LED g121 (w21) @(371,-305) /sn:0 /w:[ 3 ] /type:1
  //: LED g110 (w65) @(1472,-354) /sn:0 /w:[ 7 ] /type:1
  //: joint g60 (w55) @(611, 585) /w:[ 6 -1 12 5 ]
  _GGOR10 #(22) g29 (.I0(w40), .I1(w38), .I2(w30), .I3(w36), .I4(w35), .I5(w34), .I6(w33), .I7(w32), .I8(w56), .I9(w57), .Z(w71));   //: @(367,855) /sn:0 /w:[ 9 3 11 13 0 0 0 0 11 0 0 ]
  //: LED g168 (w29) @(-128,-114) /sn:0 /w:[ 17 ] /type:1
  _GGMUX2x8 #(8, 8) MUXPC (.I0(w15), .I1(w75), .S(w77), .Z(w0));   //: @(86,-635) /R:1 /w:[ 3 1 1 0 ] /ss:0 /do:0
  _GGMUX2x8 #(8, 8) MUXA (.I0(w9), .I1(w15), .S(w55), .Z(w4));   //: @(746,585) /w:[ 5 21 9 0 ] /ss:0 /do:0
  _GGOR11 #(24) g18 (.I0(w41), .I1(w40), .I2(w39), .I3(w30), .I4(w36), .I5(w35), .I6(w34), .I7(w33), .I8(w32), .I9(w56), .I10(w57), .Z(w7));   //: @(392,301) /sn:0 /w:[ 5 0 3 7 0 5 5 5 5 7 5 0 ]
  //: joint g199 (w15) @(276, -209) /w:[ 12 14 11 -1 ]
  //: joint g82 (w13) @(736, 363) /w:[ -1 6 8 5 ]
  demux g94 (.D0(w55), .D1(w25), .RY(w3), .PC(w75), .RF(w85));   //: @(674, 1226) /sz:(112, 102) /sn:0 /p:[ Ti0>3 Ti1>0 Ri0>5 Lo0<0 Lo1<0 ]
  //: joint g119 (w28) @(236, -394) /w:[ 2 4 -1 1 ]
  //: joint g173 (w40) @(-62, 191) /w:[ 3 4 6 -1 ]
  //: joint g107 (w59) @(832, -320) /w:[ 2 1 -1 4 ]
  //: LED g166 (w73) @(989,-62) /sn:0 /w:[ 7 ] /type:0
  //: LED g154 (w55) @(569,1031) /sn:0 /w:[ 0 ] /type:0
  //: LED g184 (w34) @(-68,419) /sn:0 /w:[ 11 ] /type:0
  //: LED g172 (w41) @(-64,137) /sn:0 /w:[ 9 ] /type:0
  //: joint g50 (w55) @(634, 585) /w:[ 8 -1 7 10 ]
  //: LED g193 (w7) @(714,65) /sn:0 /w:[ 9 ] /type:0
  //: joint g68 (w56) @(-68, 535) /w:[ 2 1 12 -1 ]
  _GGBUFIF8 #(4, 6) g9 (.Z(w65), .I(w48), .E(w73));   //: @(1485,851) /sn:0 /w:[ 0 5 13 ]
  //: joint g73 (w73) @(1091, 744) /w:[ 10 9 16 -1 ]
  //: LED g133 (w10) @(615,-258) /sn:0 /w:[ 3 ] /type:1
  _GGMUX2x8 #(8, 8) MUXB (.I0(w37), .I1(w60), .S(w55), .Z(w5));   //: @(933,585) /w:[ 5 0 11 0 ] /ss:0 /do:0
  //: joint g59 (w55) @(611, 1054) /w:[ 2 4 1 -1 ]
  //: joint g102 (w69) @(1026, 860) /w:[ 2 12 -1 1 ]
  //: joint g22 (w56) @(160, 535) /w:[ 6 -1 5 8 ]
  //: joint g31 (w56) @(52, 535) /w:[ 4 -1 3 10 ]
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g71 (.A(w62), .D(w48), .WE(w73), .OE(w69), .CS(~w78));   //: @(1243,787) /sn:0 /w:[ 0 0 15 9 1 ]
  //: joint g169 (w29) @(-128, -49) /w:[ 2 16 1 -1 ]
  //: LED g186 (w33) @(-69,452) /sn:0 /w:[ 11 ] /type:0
  //: LED g87 (w60) @(988,538) /sn:0 /w:[ 3 ] /type:1
  //: LED g99 (w73) @(1023,723) /sn:0 /w:[ 23 ] /type:0
  //: LED g83 (w37) @(1021,470) /sn:0 /w:[ 3 ] /type:1
  _GGOR4 #(10) g203 (.I0(w44), .I1(w43), .I2(w81), .I3(w45), .Z(w77));   //: @(-86,-272) /sn:0 /R:1 /w:[ 3 0 0 0 0 ]
  //: joint g36 (w36) @(23, 361) /w:[ 1 -1 2 12 ]
  //: SWITCH g41 (w52) @(644,454) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g45 (w53) @(643,394) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g69 (w32) @(-69, 506) /w:[ 9 10 12 -1 ]
  //: joint g213 (w73) @(1243, 744) /w:[ 12 -1 11 14 ]
  //: joint g42 (w52) @(679, 454) /w:[ 2 4 1 -1 ]
  //: LED g138 (w81) @(-5,50) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: LED g156 (w25) @(815,1029) /sn:0 /w:[ 3 ] /type:0
  //: LED g66 (w14) @(970,329) /sn:0 /w:[ 3 ] /type:1
  //: LED g151 (w4) @(1375,495) /sn:0 /w:[ 3 ] /type:1
  //: joint g167 (w73) @(989, -33) /w:[ 4 6 3 -1 ]
  //: joint g153 (w15) @(236, -267) /w:[ -1 1 2 4 ]
  //: joint g146 (w5) @(933, 672) /w:[ 2 1 -1 4 ]
  //: LED g162 (w7) @(441,268) /sn:0 /w:[ 11 ] /type:0
  //: LED g191 (w57) @(-67,548) /sn:0 /w:[ 11 ] /type:0
  //: joint g28 (w41) @(61, 157) /w:[ 4 -1 3 6 ]
  //: joint g34 (w34) @(34, 441) /w:[ 2 -1 8 1 ]
  //: joint g46 (w53) @(790, 394) /w:[ 2 -1 1 4 ]
  //: SWITCH g57 (w54) @(969,947) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: GROUND g118 (w27) @(299,-511) /sn:0 /R:1 /w:[ 1 ]
  //: joint g84 (w37) @(923, 493) /w:[ 2 1 -1 4 ]
  //: SWITCH g5 (w18) @(637,-323) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g11 (w24) @(685,258) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGMUX2x3 #(8, 8) g14 (.I0(w11), .I1(w10), .S(w73), .Z(w12));   //: @(1027,34) /sn:0 /R:3 /w:[ 0 0 5 3 ] /ss:0 /do:0
  //: joint g150 (w62) @(1190, 788) /w:[ 1 2 4 -1 ]
  //: joint g112 (w4) @(746, 634) /w:[ 2 1 -1 4 ]
  //: SWITCH g201 (w50) @(407,-116) /sn:0 /w:[ 1 ] /st:1 /dn:1
  //: LED g123 (w1) @(637,-89) /sn:0 /w:[ 3 ] /type:1
  _GGAND3 #(8) g61 (.I0(w7), .I1(w71), .I2(w76), .Z(w68));   //: @(441,973) /sn:0 /w:[ 13 13 1 0 ]
  //: joint g21 (w57) @(152, 564) /w:[ 4 -1 3 6 ]
  //: LED g187 (w32) @(-69,486) /sn:0 /w:[ 11 ] /type:0
  //: LED g115 (w28) @(331,-409) /sn:0 /w:[ 3 ] /type:1
  _GGOR8 #(18) g20 (.I0(w41), .I1(w30), .I2(w35), .I3(w34), .I4(w33), .I5(w32), .I6(w56), .I7(w57), .Z(w64));   //: @(390,578) /sn:0 /w:[ 7 9 7 7 7 7 9 7 0 ]
  //: joint g32 (w32) @(46, 506) /w:[ 2 -1 8 1 ]
  //: LED g79 (w49) @(971,799) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g97 (w36) @(-65, 361) /w:[ 5 6 8 -1 ]
  //: joint g134 (w10) @(615, -138) /w:[ 1 2 4 -1 ]
  //: LED g145 (w5) @(1004,652) /sn:0 /w:[ 3 ] /type:1
  //: LED g175 (w39) @(-66,203) /sn:0 /w:[ 5 ] /type:0
  //: joint g148 (w69) @(1250, 833) /w:[ 6 8 -1 5 ]
  //: LED g89 (w15) @(671,536) /sn:0 /w:[ 19 ] /type:1
  dec_4to16 g15 (.a(w29), .y15(w45), .y14(w81), .y13(w43), .y12(w44), .y11(w41), .y10(w40), .y9(w39), .y8(w38), .y7(w30), .y6(w36), .y5(w35), .y4(w34), .y3(w33), .y2(w32), .y1(w56), .y0(w57));   //: @(-265, -9) /sz:(189, 590) /sn:0 /p:[ Li0>0 Ro0<5 Ro1<5 Ro2<5 Ro3<5 Ro4<0 Ro5<7 Ro6<0 Ro7<0 Ro8<0 Ro9<9 Ro10<13 Ro11<13 Ro12<13 Ro13<13 Ro14<13 Ro15<13 ]
  //: LED g129 (w62) @(968,-282) /sn:0 /w:[ 7 ] /type:1
  //: joint g147 (w38) @(-68, 271) /w:[ 2 4 1 -1 ]
  //: joint g27 (w30) @(84, 312) /w:[ 6 -1 5 8 ]
  //: joint g165 (w12) @(938, 34) /w:[ 2 4 1 -1 ]
  //: joint g62 (w3) @(831, 1042) /w:[ 2 1 -1 4 ]
  //: LED g160 (w64) @(453,552) /sn:0 /w:[ 9 ] /type:0
  //: joint g171 (w0) @(223, -671) /w:[ 2 4 1 -1 ]
  //: joint g88 (w60) @(943, 556) /w:[ 2 4 -1 1 ]
  //: joint g55 (w29) @(429, 41) /w:[ 4 -1 3 10 ]
  //: LED g195 (w64) @(677,65) /sn:0 /w:[ 7 ] /type:0
  assign w2 = w16[8:6]; //: TAP g13 @(515,15) /sn:0 /R:2 /w:[ 5 18 17 ] /ss:1
  assign w55 = w16[2]; //: TAP g53 @(515,-54) /sn:0 /R:2 /w:[ 13 14 13 ] /ss:0
  //: LED g135 (w29) @(445,-31) /sn:0 /w:[ 9 ] /type:1
  //: LED g139 (w43) @(-3,81) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: LED g140 (w44) @(-3,117) /sn:0 /R:3 /w:[ 0 ] /type:0

endmodule
//: /netlistEnd

//: /netlistBegin final_sub
module final_sub(S, B, A, COUT);
//: interface  /sz:(117, 103) /bd:[ Li0>B[7:0](68/103) Li1>A[7:0](34/103) Ro0<S[7:0](68/103) Ro1<COUT(34/103) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:603,295)(460,295)(460,295)(450,295){1}
//: {2}(448,293)(448,235)(448,235)(448,163){3}
//: {4}(450,161)(#:602,161){5}
//: {6}(448,159)(448,113){7}
//: {8}(448,297)(448,303)(448,303)(#:448,375){9}
output COUT;    //: /sn:0 {0}(698,267)(837,267)(837,259)(847,259){1}
//: {2}(851,259)(861,259)(861,259)(910,259){3}
//: {4}(849,257)(849,251){5}
//: {6}(849,261)(849,268){7}
input [7:0] A;    //: /sn:0 {0}(#:603,267)(417,267)(417,267)(413,267){1}
//: {2}(411,265)(411,233)(411,233)(411,191){3}
//: {4}(413,189)(#:602,189){5}
//: {6}(411,187)(411,108){7}
//: {8}(411,269)(411,286)(411,286)(#:411,372){9}
output [7:0] S;    //: /sn:0 {0}(#:862,228)(888,228)(888,228)(903,228){1}
wire w4;    //: /sn:0 {0}(697,161)(761,161)(761,108)(771,108){1}
//: {2}(775,108)(822,108)(822,107){3}
//: {4}(773,110)(773,115){5}
wire [7:0] w1;    //: /sn:0 {0}(#:697,189)(809,189)(809,218)(833,218){1}
wire [7:0] w2;    //: /sn:0 {0}(#:698,295)(818,295)(818,238)(833,238){1}
//: enddecls

  sub_8 g8 (.A(B), .B(A), .cout(w4), .s(w1));   //: @(603, 134) /sz:(93, 83) /sn:0 /p:[ Li0>5 Li1>5 Ro0<0 Ro1<0 ]
  //: OUT g4 (S) @(900,228) /sn:0 /w:[ 1 ]
  //: IN g3 (B) @(448,377) /sn:0 /R:1 /w:[ 9 ]
  //: IN g2 (A) @(411,374) /sn:0 /R:1 /w:[ 9 ]
  //: joint g1 (COUT) @(849, 259) /w:[ 2 4 1 6 ]
  //: joint g10 (B) @(448, 161) /w:[ 4 6 -1 3 ]
  //: LED g6 (w4) @(822,100) /sn:0 /w:[ 3 ] /type:0
  sub_8 g9 (.A(A), .B(B), .cout(COUT), .s(w2));   //: @(604, 240) /sz:(93, 83) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<0 ]
  //: joint g7 (w4) @(773, 108) /w:[ 2 -1 1 4 ]
  //: joint g12 (A) @(411, 267) /w:[ 1 2 -1 8 ]
  //: joint g11 (A) @(411, 189) /w:[ 4 6 -1 3 ]
  //: OUT g5 (COUT) @(907,259) /sn:0 /w:[ 3 ]
  _GGMUX2x8 #(8, 8) g0 (.I0(w2), .I1(w1), .S(COUT), .Z(S));   //: @(849,228) /sn:0 /R:1 /w:[ 1 1 5 0 ] /ss:0 /do:0
  //: joint g13 (B) @(448, 295) /w:[ 1 2 -1 8 ]

endmodule
//: /netlistEnd

//: /netlistBegin dec
module dec(w9, w4, w5, w22, w7, w1, w8, w0, w26, w20, w3, w6, w10, w25, w23, w24, w2, w21);
//: interface  /sz:(291, 259) /bd:[ Li0>w10(30/259) Li1>w1[2:0](15/259) Ro0<w26(243/259) Ro1<w25(228/259) Ro2<w24(213/259) Ro3<w23(198/259) Ro4<w22(182/259) Ro5<w21(167/259) Ro6<w20(152/259) Ro7<w9(137/259) Ro8<w8(121/259) Ro9<w7(106/259) Ro10<w6(91/259) Ro11<w5(76/259) Ro12<w4(60/259) Ro13<w3(45/259) Ro14<w2(30/259) Ro15<w0(15/259) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output w6;    //: /sn:0 {0}(480,378)(407,378)(407,379)(366,379){1}
output w7;    //: /sn:0 {0}(424,375)(381,375)(381,372)(366,372){1}
output w25;    //: /sn:0 {0}(364,501)(462,501){1}
output w4;    //: /sn:0 {0}(488,494)(364,494){1}
output w22;    //: /sn:0 {0}(364,508)(483,508)(483,507)(498,507){1}
output w3;    //: /sn:0 {0}(431,415)(381,415)(381,399)(366,399){1}
output w0;    //: /sn:0 {0}(423,349)(381,349)(381,352)(366,352){1}
output w20;    //: /sn:0 {0}(417,396)(381,396)(381,392)(366,392){1}
output w23;    //: /sn:0 {0}(364,521)(392,521)(392,519)(407,519){1}
input w10;    //: /sn:0 {0}(188,410)(300,410)(300,413){1}
//: {2}(302,415)(350,415)(350,398){3}
//: {4}(300,417)(300,425)(301,425)(301,434){5}
output w24;    //: /sn:0 {0}(364,528)(403,528)(403,533)(418,533){1}
output w21;    //: /sn:0 {0}(473,387)(418,387)(418,385)(366,385){1}
input [2:0] w1;    //: /sn:0 {0}(#:183,371)(203,371)(203,376)(255,376){1}
//: {2}(259,376)(337,376){3}
//: {4}(#:257,378)(257,505)(335,505){5}
output w8;    //: /sn:0 {0}(444,368)(412,368)(412,365)(366,365){1}
output w2;    //: /sn:0 {0}(467,481)(364,481){1}
output w5;    //: /sn:0 {0}(364,488)(396,488){1}
output w26;    //: /sn:0 {0}(364,514)(456,514)(456,515)(471,515){1}
output w9;    //: /sn:0 {0}(431,360)(381,360)(381,359)(366,359){1}
wire w11;    //: /sn:0 {0}(301,450)(301,542)(348,542)(348,527){1}
//: enddecls

  //: OUT g8 (w9) @(428,360) /sn:0 /w:[ 0 ]
  //: joint g4 (w1) @(257, 376) /w:[ 2 -1 1 4 ]
  //: OUT g16 (w4) @(485,494) /sn:0 /w:[ 0 ]
  //: joint g3 (w10) @(300, 415) /w:[ 2 1 -1 4 ]
  //: OUT g17 (w5) @(393,488) /sn:0 /w:[ 1 ]
  _GGNBUF #(2) g2 (.I(w10), .Z(w11));   //: @(301,440) /sn:0 /R:3 /w:[ 5 0 ]
  _GGDECODER8 #(6, 6) g1 (.I(w1), .E(w11), .Z0(w24), .Z1(w23), .Z2(w26), .Z3(w22), .Z4(w25), .Z5(w4), .Z6(w5), .Z7(w2));   //: @(348,505) /sn:0 /R:1 /w:[ 5 1 0 0 0 0 0 1 0 1 ] /ss:0 /do:0
  //: OUT g18 (w22) @(495,507) /sn:0 /w:[ 1 ]
  //: OUT g10 (w7) @(421,375) /sn:0 /w:[ 0 ]
  //: IN g6 (w1) @(181,371) /sn:0 /w:[ 0 ]
  //: OUT g9 (w8) @(441,368) /sn:0 /w:[ 0 ]
  //: OUT g7 (w0) @(420,349) /sn:0 /w:[ 0 ]
  //: OUT g22 (w26) @(468,515) /sn:0 /w:[ 1 ]
  //: OUT g12 (w20) @(414,396) /sn:0 /w:[ 0 ]
  //: OUT g14 (w3) @(428,415) /sn:0 /w:[ 0 ]
  //: OUT g11 (w6) @(477,378) /sn:0 /w:[ 0 ]
  //: IN g5 (w10) @(186,410) /sn:0 /w:[ 0 ]
  //: OUT g21 (w25) @(459,501) /sn:0 /w:[ 1 ]
  //: OUT g19 (w23) @(404,519) /sn:0 /w:[ 1 ]
  //: OUT g20 (w24) @(415,533) /sn:0 /w:[ 1 ]
  //: OUT g15 (w2) @(464,481) /sn:0 /w:[ 0 ]
  _GGDECODER8 #(6, 6) g0 (.I(w1), .E(w10), .Z0(w3), .Z1(w20), .Z2(w21), .Z3(w6), .Z4(w7), .Z5(w8), .Z6(w9), .Z7(w0));   //: @(350,376) /sn:0 /R:1 /w:[ 3 3 1 1 1 1 1 1 1 1 ] /ss:0 /do:0
  //: OUT g13 (w21) @(470,387) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin comp4
module comp4(b1, b2, g, b3, a1, l, e, a0, a2, a3, b0);
//: interface  /sz:(111, 261) /bd:[ Li0>a0(29/261) Li1>a1(58/261) Li2>a2(87/261) Li3>a3(116/261) Li4>b0(145/261) Li5>b1(174/261) Li6>b2(203/261) Li7>b3(232/261) Ro0<e(29/261) Ro1<g(58/261) Ro2<l(87/261) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(-247,614)(-170,614){1}
//: {2}(-166,614)(-144,614){3}
//: {4}(-168,616)(-168,662)(-86,662){5}
input b2;    //: /sn:0 {0}(-245,667)(-179,667){1}
//: {2}(-175,667)(-144,667){3}
//: {4}(-177,665)(-177,619)(-86,619){5}
input a3;    //: /sn:0 {0}(-248,510)(-173,510){1}
//: {2}(-169,510)(-144,510){3}
//: {4}(-171,512)(-171,553)(-87,553){5}
output l;    //: /sn:0 {0}(282,693)(249,693)(249,693)(342,693){1}
input b3;    //: /sn:0 {0}(-249,558)(-181,558){1}
//: {2}(-177,558)(-144,558){3}
//: {4}(-179,556)(-179,515)(-86,515){5}
input a1;    //: /sn:0 {0}(-242,722)(-168,722){1}
//: {2}(-164,722)(-144,722){3}
//: {4}(-166,724)(-166,771)(-86,771){5}
input b1;    //: /sn:0 {0}(-242,776)(-177,776){1}
//: {2}(-173,776)(-144,776){3}
//: {4}(-175,774)(-175,727)(-86,727){5}
input a0;    //: /sn:0 {0}(-86,872)(-164,872)(-164,823){1}
//: {2}(-162,821)(-144,821){3}
//: {4}(-166,821)(-241,821){5}
input b0;    //: /sn:0 {0}(-239,877)(-176,877){1}
//: {2}(-172,877)(-144,877){3}
//: {4}(-174,875)(-174,826)(-86,826){5}
output e;    //: /sn:0 {0}(127,933)(309,933)(309,933)(347,933){1}
output g;    //: /sn:0 {0}(279,837)(298,837)(298,837)(344,837){1}
wire w16;    //: /sn:0 {0}(-65,617)(-16,617){1}
//: {2}(-14,615)(-14,577)(106,577){3}
//: {4}(-14,619)(-14,636)(1,636){5}
wire w6;    //: /sn:0 {0}(106,931)(58,931)(58,877){1}
//: {2}(60,875)(106,875){3}
//: {4}(58,873)(58,823){5}
//: {6}(60,821)(106,821){7}
//: {8}(58,819)(58,769){9}
//: {10}(60,767)(106,767){11}
//: {12}(58,765)(58,715){13}
//: {14}(60,713)(106,713){15}
//: {16}(58,711)(58,639)(22,639){17}
wire w7;    //: /sn:0 {0}(-128,667)(-86,667){1}
wire w34;    //: /sn:0 {0}(258,840)(217,840)(217,767)(127,767){1}
wire w25;    //: /sn:0 {0}(106,772)(48,772)(48,774)(-11,774){1}
//: {2}(-13,772)(-13,750)(1,750){3}
//: {4}(-15,774)(-65,774){5}
wire w4;    //: /sn:0 {0}(-65,513)(-16,513){1}
//: {2}(-12,513)(253,513)(253,686)(261,686){3}
//: {4}(-14,515)(-14,531)(1,531){5}
wire w3;    //: /sn:0 {0}(-128,558)(-87,558){1}
wire w22;    //: /sn:0 {0}(106,718)(-14,718)(-14,723){1}
//: {2}(-16,725)(-65,725){3}
//: {4}(-14,727)(-14,745)(1,745){5}
wire w0;    //: /sn:0 {0}(106,926)(65,926)(65,872){1}
//: {2}(67,870)(106,870){3}
//: {4}(65,868)(65,818){5}
//: {6}(67,816)(106,816){7}
//: {8}(65,814)(65,764){9}
//: {10}(67,762)(106,762){11}
//: {12}(65,760)(65,710){13}
//: {14}(67,708)(106,708){15}
//: {16}(65,706)(65,662){17}
//: {18}(67,660)(106,660){19}
//: {20}(65,658)(65,574){21}
//: {22}(67,572)(106,572){23}
//: {24}(65,570)(65,534)(22,534){25}
wire w30;    //: /sn:0 {0}(-128,877)(-86,877){1}
wire w37;    //: /sn:0 {0}(127,713)(246,713)(246,696)(261,696){1}
wire w19;    //: /sn:0 {0}(-65,665)(-16,665){1}
//: {2}(-12,665)(106,665){3}
//: {4}(-14,663)(-14,641)(1,641){5}
wire w23;    //: /sn:0 {0}(127,877)(243,877)(243,845)(258,845){1}
wire w10;    //: /sn:0 {0}(-66,556)(-16,556){1}
//: {2}(-12,556)(233,556)(233,830)(258,830){3}
//: {4}(-14,554)(-14,536)(1,536){5}
wire w24;    //: /sn:0 {0}(-128,776)(-86,776){1}
wire w31;    //: /sn:0 {0}(106,885)(-15,885)(-15,877){1}
//: {2}(-15,873)(-15,852)(0,852){3}
//: {4}(-17,875)(-65,875){5}
wire w1;    //: /sn:0 {0}(-128,510)(-86,510){1}
wire w8;    //: /sn:0 {0}(127,575)(246,575)(246,691)(261,691){1}
wire w17;    //: /sn:0 {0}(106,936)(51,936)(51,882){1}
//: {2}(53,880)(106,880){3}
//: {4}(51,878)(51,828){5}
//: {6}(53,826)(106,826){7}
//: {8}(51,824)(51,748)(22,748){9}
wire w28;    //: /sn:0 {0}(106,831)(-13,831){1}
//: {2}(-15,829)(-15,824)(-65,824){3}
//: {4}(-15,833)(-15,847)(0,847){5}
wire w11;    //: /sn:0 {0}(-128,821)(-86,821){1}
wire w2;    //: /sn:0 {0}(127,823)(251,823)(251,701)(261,701){1}
wire w15;    //: /sn:0 {0}(-128,722)(-86,722){1}
wire w5;    //: /sn:0 {0}(-128,614)(-86,614){1}
wire w9;    //: /sn:0 {0}(21,850)(45,850)(45,941)(106,941){1}
wire w40;    //: /sn:0 {0}(127,663)(224,663)(224,835)(258,835){1}
//: enddecls

  _GGNBUF #(2) g4 (.I(b1), .Z(w24));   //: @(-138,776) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g8 (.I0(w1), .I1(b3), .Z(w4));   //: @(-75,513) /sn:0 /w:[ 1 5 0 ]
  _GGAND3 #(8) g44 (.I0(w0), .I1(w6), .I2(w22), .Z(w37));   //: @(117,713) /sn:0 /w:[ 15 15 0 0 ]
  //: IN g16 (b1) @(-244,776) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g3 (.I(b2), .Z(w7));   //: @(-138,667) /sn:0 /w:[ 3 0 ]
  //: joint g47 (w0) @(65, 816) /w:[ 6 8 -1 5 ]
  //: IN g17 (b2) @(-247,667) /sn:0 /w:[ 0 ]
  //: joint g26 (b2) @(-177, 667) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g2 (.I(a2), .Z(w5));   //: @(-138,614) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g23 (.I0(a0), .I1(w30), .Z(w31));   //: @(-75,875) /sn:0 /w:[ 0 1 5 ]
  //: joint g30 (a1) @(-166, 722) /w:[ 2 -1 1 4 ]
  //: OUT g39 (g) @(341,837) /sn:0 /w:[ 1 ]
  _GGNBUF #(2) g1 (.I(b3), .Z(w3));   //: @(-138,558) /sn:0 /w:[ 3 0 ]
  //: joint g24 (b3) @(-179, 558) /w:[ 2 4 1 -1 ]
  //: joint g29 (b1) @(-175, 776) /w:[ 2 4 1 -1 ]
  //: joint g60 (w6) @(58, 875) /w:[ 2 4 -1 1 ]
  //: joint g51 (w0) @(65, 572) /w:[ 22 24 -1 21 ]
  //: IN g18 (b3) @(-251,558) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g10 (.I0(w5), .I1(b2), .Z(w16));   //: @(-75,617) /sn:0 /w:[ 1 5 0 ]
  //: joint g25 (a3) @(-171, 510) /w:[ 2 -1 1 4 ]
  _GGOR4 #(10) g65 (.I0(w10), .I1(w40), .I2(w34), .I3(w23), .Z(g));   //: @(269,837) /sn:0 /w:[ 3 1 0 1 0 ]
  _GGOR4 #(10) g64 (.I0(w4), .I1(w8), .I2(w37), .I3(w2), .Z(l));   //: @(272,693) /sn:0 /w:[ 3 1 1 1 0 ]
  //: joint g49 (w0) @(65, 708) /w:[ 14 16 -1 13 ]
  _GGNBUF #(2) g6 (.I(b0), .Z(w30));   //: @(-138,877) /sn:0 /w:[ 3 0 ]
  //: joint g50 (w0) @(65, 762) /w:[ 10 12 -1 9 ]
  _GGNBUF #(2) g7 (.I(a1), .Z(w15));   //: @(-138,722) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g9 (.I0(a3), .I1(w3), .Z(w10));   //: @(-76,556) /sn:0 /w:[ 5 1 0 ]
  _GGNOR2 #(4) g35 (.I0(w28), .I1(w31), .Z(w9));   //: @(11,850) /sn:0 /w:[ 5 3 0 ]
  //: joint g56 (w25) @(-13, 774) /w:[ 1 2 4 -1 ]
  //: joint g58 (w28) @(-15, 831) /w:[ 1 2 -1 4 ]
  //: IN g22 (a1) @(-244,722) /sn:0 /w:[ 0 ]
  //: joint g31 (b0) @(-174, 877) /w:[ 2 4 1 -1 ]
  //: joint g59 (w31) @(-15, 875) /w:[ -1 2 4 1 ]
  //: joint g67 (w10) @(-14, 556) /w:[ 2 4 1 -1 ]
  //: OUT g41 (l) @(339,693) /sn:0 /w:[ 1 ]
  _GGNOR2 #(4) g33 (.I0(w16), .I1(w19), .Z(w6));   //: @(12,639) /sn:0 /w:[ 5 5 17 ]
  _GGAND2 #(6) g36 (.I0(w0), .I1(w16), .Z(w8));   //: @(117,575) /sn:0 /w:[ 23 3 0 ]
  _GGAND2 #(6) g45 (.I0(w0), .I1(w19), .Z(w40));   //: @(117,663) /sn:0 /w:[ 19 3 0 ]
  //: joint g54 (w6) @(58, 713) /w:[ 14 16 -1 13 ]
  //: OUT g40 (e) @(344,933) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g42 (.I0(w0), .I1(w6), .I2(w17), .I3(w28), .Z(w2));   //: @(117,823) /sn:0 /w:[ 7 7 7 0 0 ]
  //: joint g52 (w16) @(-14, 617) /w:[ -1 2 1 4 ]
  //: joint g66 (w4) @(-14, 513) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g12 (.I0(w15), .I1(b1), .Z(w22));   //: @(-75,725) /sn:0 /w:[ 1 5 3 ]
  //: joint g28 (a0) @(-164, 821) /w:[ 2 -1 4 1 ]
  _GGNOR2 #(4) g34 (.I0(w22), .I1(w25), .Z(w17));   //: @(12,748) /sn:0 /w:[ 5 3 9 ]
  //: joint g46 (w0) @(65, 870) /w:[ 2 4 -1 1 ]
  //: joint g57 (w6) @(58, 767) /w:[ 10 12 -1 9 ]
  //: IN g14 (a0) @(-243,821) /sn:0 /w:[ 5 ]
  _GGNBUF #(2) g5 (.I(a0), .Z(w11));   //: @(-138,821) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g11 (.I0(a2), .I1(w7), .Z(w19));   //: @(-75,665) /sn:0 /w:[ 5 1 0 ]
  //: IN g19 (a2) @(-249,614) /sn:0 /w:[ 0 ]
  //: IN g21 (a3) @(-250,510) /sn:0 /w:[ 0 ]
  //: joint g61 (w17) @(51, 880) /w:[ 2 4 -1 1 ]
  //: IN g20 (b0) @(-241,877) /sn:0 /w:[ 0 ]
  _GGNOR2 #(4) g32 (.I0(w4), .I1(w10), .Z(w0));   //: @(12,534) /sn:0 /w:[ 5 5 25 ]
  //: joint g63 (w17) @(51, 826) /w:[ 6 8 -1 5 ]
  _GGNBUF #(2) g0 (.I(a3), .Z(w1));   //: @(-138,510) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g15 (.I0(w11), .I1(b0), .Z(w28));   //: @(-75,824) /sn:0 /w:[ 1 5 3 ]
  _GGAND4 #(10) g38 (.I0(w0), .I1(w6), .I2(w17), .I3(w31), .Z(w23));   //: @(117,877) /sn:0 /w:[ 3 3 3 0 0 ]
  _GGAND3 #(8) g43 (.I0(w0), .I1(w6), .I2(w25), .Z(w34));   //: @(117,767) /sn:0 /w:[ 11 11 0 1 ]
  //: joint g27 (a2) @(-168, 614) /w:[ 2 -1 1 4 ]
  //: joint g48 (w0) @(65, 660) /w:[ 18 20 -1 17 ]
  _GGAND4 #(10) g37 (.I0(w0), .I1(w6), .I2(w17), .I3(w9), .Z(e));   //: @(117,933) /sn:0 /w:[ 0 0 0 1 0 ]
  //: joint g62 (w6) @(58, 821) /w:[ 6 8 -1 5 ]
  //: joint g55 (w22) @(-14, 725) /w:[ -1 1 2 4 ]
  _GGAND2 #(6) g13 (.I0(a1), .I1(w24), .Z(w25));   //: @(-75,774) /sn:0 /w:[ 5 1 5 ]
  //: joint g53 (w19) @(-14, 665) /w:[ 2 4 1 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin comp
module comp(b, a, et, lt, gt);
//: interface  /sz:(148, 189) /bd:[ Li0>a[7:0](47/189) Li1>b[7:0](94/189) Ro0<et(86/189) Ro1<gt(34/189) Ro2<lt(141/189) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output et;    //: /sn:0 {0}(640,121)(722,121)(722,117)(737,117){1}
input [7:0] b;    //: /sn:0 {0}(#:-4,507)(-4,489){1}
//: {2}(-4,488)(-4,443){3}
//: {4}(-4,442)(-4,402){5}
//: {6}(-4,401)(-4,358){7}
//: {8}(-4,357)(-4,69){9}
//: {10}(-4,68)(-4,23){11}
//: {12}(-4,22)(-4,-18){13}
//: {14}(-4,-19)(-4,-62){15}
//: {16}(-4,-63)(-4,-283){17}
output lt;    //: /sn:0 {0}(640,407)(737,407){1}
input [7:0] a;    //: /sn:0 {0}(#:-66,513)(-66,287){1}
//: {2}(-66,286)(-66,249){3}
//: {4}(-66,248)(-66,206){5}
//: {6}(-66,205)(-66,185)(-65,185)(-65,163){7}
//: {8}(-65,162)(-65,15)(-66,15)(-66,-133){9}
//: {10}(-66,-134)(-66,-171){11}
//: {12}(-66,-172)(-66,-214){13}
//: {14}(-66,-215)(-66,-258){15}
//: {16}(-66,-259)(-66,-285){17}
output gt;    //: /sn:0 {0}(640,-167)(722,-167)(722,-169)(737,-169){1}
wire w16;    //: /sn:0 {0}(-62,206)(127,206)(127,524)(163,524){1}
wire w13;    //: /sn:0 {0}(0,443)(120,443)(120,761)(163,761){1}
wire w6;    //: /sn:0 {0}(-62,-171)(164,-171){1}
wire w7;    //: /sn:0 {0}(-62,-133)(164,-133){1}
wire w4;    //: /sn:0 {0}(-62,-258)(164,-258){1}
wire w25;    //: /sn:0 {0}(544,319)(604,319)(604,404)(619,404){1}
wire w0;    //: /sn:0 {0}(0,-62)(164,-62){1}
wire w3;    //: /sn:0 {0}(0,69)(164,69){1}
wire w20;    //: /sn:0 {0}(495,-113)(485,-113)(485,-98)(514,-98)(514,551)(315,551){1}
wire w18;    //: /sn:0 {0}(-62,287)(211,287)(211,300){1}
//: {2}(209,302)(203,302){3}
//: {4}(211,304)(211,314)(153,314)(153,605)(163,605){5}
wire w12;    //: /sn:0 {0}(209,417)(214,417){1}
//: {2}(216,415)(216,402)(0,402){3}
//: {4}(216,419)(216,429)(155,429)(155,720)(163,720){5}
wire w19;    //: /sn:0 {0}(523,321)(513,321)(513,336)(532,336)(532,885)(362,885)(362,726)(332,726)(332,714)(315,714){1}
wire w10;    //: /sn:0 {0}(619,118)(518,118){1}
//: {2}(514,118)(403,118)(403,-115){3}
//: {4}(405,-117)(415,-117)(415,-118)(495,-118){5}
//: {6}(401,-117)(357,-117)(357,-113)(316,-113){7}
//: {8}(516,120)(516,316)(523,316){9}
wire w23;    //: /sn:0 {0}(516,-115)(604,-115)(604,-165)(619,-165){1}
wire w21;    //: /sn:0 {0}(619,123)(609,123)(609,138)(641,138)(641,724)(355,724)(355,625)(315,625){1}
wire w1;    //: /sn:0 {0}(0,-18)(164,-18){1}
wire w8;    //: /sn:0 {0}(619,409)(441,409)(441,-24)(316,-24){1}
wire w17;    //: /sn:0 {0}(-62,249)(142,249)(142,567)(163,567){1}
wire w14;    //: /sn:0 {0}(0,489)(131,489)(131,807)(163,807){1}
wire w11;    //: /sn:0 {0}(0,358)(216,358)(216,371){1}
//: {2}(214,373)(208,373){3}
//: {4}(216,375)(216,385)(155,385)(155,676)(163,676){5}
wire w2;    //: /sn:0 {0}(0,23)(164,23){1}
wire w15;    //: /sn:0 {0}(-70,163)(-104,163)(-104,480)(163,480){1}
wire w5;    //: /sn:0 {0}(-62,-214)(164,-214){1}
wire w9;    //: /sn:0 {0}(316,-187)(602,-187)(602,-170)(619,-170){1}
//: enddecls

  assign w14 = b[0]; //: TAP g4 @(-6,489) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  assign w15 = a[3]; //: TAP g8 @(-67,163) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:0
  //: IN g3 (b) @(-4,509) /sn:0 /R:1 /w:[ 0 ]
  assign w4 = a[7]; //: TAP g16 @(-68,-258) /sn:0 /R:2 /w:[ 0 15 16 ] /ss:1
  assign w7 = a[4]; //: TAP g17 @(-68,-133) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1
  //: joint g26 (w10) @(516, 118) /w:[ 1 -1 2 8 ]
  //: IN g2 (a) @(-66,515) /sn:0 /R:1 /w:[ 0 ]
  _GGAND2 #(6) g23 (.I0(w10), .I1(w20), .Z(w23));   //: @(506,-115) /sn:0 /w:[ 5 0 0 ]
  comp4 g30 (.a0(w18), .a1(w17), .a2(w16), .a3(w15), .b0(w14), .b1(w13), .b2(w12), .b3(w11), .e(w21), .g(w20), .l(w19));   //: @(164, 426) /sz:(150, 410) /sn:0 /p:[ Li0>5 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>5 Li7>5 Ro0<1 Ro1<1 Ro2<1 ]
  _GGAND2 #(6) g24 (.I0(w10), .I1(w19), .Z(w25));   //: @(534,319) /sn:0 /w:[ 9 0 0 ]
  //: joint g1 (w18) @(211, 302) /w:[ -1 1 2 4 ]
  //: OUT g29 (et) @(734,117) /sn:0 /w:[ 1 ]
  assign w6 = a[5]; //: TAP g18 @(-68,-171) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  assign w17 = a[1]; //: TAP g10 @(-68,249) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: joint g25 (w10) @(403, -117) /w:[ 4 -1 6 3 ]
  assign w12 = b[2]; //: TAP g6 @(-6,402) /sn:0 /R:2 /w:[ 3 5 6 ] /ss:1
  assign w11 = b[3]; //: TAP g7 @(-6,358) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  assign w16 = a[2]; //: TAP g9 @(-68,206) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  _GGAND2 #(6) g22 (.I0(w10), .I1(w21), .Z(et));   //: @(630,121) /sn:0 /w:[ 0 0 0 ]
  //: joint g31 (w11) @(216, 373) /w:[ -1 1 2 4 ]
  assign w0 = b[7]; //: TAP g12 @(-6,-62) /sn:0 /R:2 /w:[ 0 15 16 ] /ss:1
  //: OUT g28 (lt) @(734,407) /sn:0 /w:[ 1 ]
  assign w13 = b[1]; //: TAP g5 @(-6,443) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  assign w18 = a[0]; //: TAP g11 @(-68,287) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  assign w2 = b[5]; //: TAP g14 @(-6,23) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  assign w5 = a[6]; //: TAP g19 @(-68,-214) /sn:0 /R:2 /w:[ 0 13 14 ] /ss:1
  _GGOR2 #(6) g21 (.I0(w25), .I1(w8), .Z(lt));   //: @(630,407) /sn:0 /w:[ 1 0 0 ]
  _GGOR2 #(6) g20 (.I0(w9), .I1(w23), .Z(gt));   //: @(630,-167) /sn:0 /w:[ 1 1 0 ]
  //: joint g32 (w12) @(216, 417) /w:[ -1 2 1 4 ]
  comp4 g0 (.a0(w7), .a1(w6), .a2(w5), .a3(w4), .b0(w3), .b1(w2), .b2(w1), .b3(w0), .e(w10), .g(w9), .l(w8));   //: @(165, -312) /sz:(150, 410) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>1 Li7>1 Ro0<7 Ro1<0 Ro2<1 ]
  assign w1 = b[6]; //: TAP g15 @(-6,-18) /sn:0 /R:2 /w:[ 0 13 14 ] /ss:1
  //: OUT g27 (gt) @(734,-169) /sn:0 /w:[ 1 ]
  assign w3 = b[4]; //: TAP g13 @(-6,69) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin dec_4to16
module dec_4to16(y4, y14, y5, a, y11, y12, y6, y13, y10, y0, y2, y9, y7, y8, y3, y15, y1);
//: interface  /sz:(189, 590) /bd:[ Li0>a[3:0](34/590) Ro0<y0(573/590) Ro1<y1(544/590) Ro2<y2(515/590) Ro3<y3(481/590) Ro4<y4(450/590) Ro5<y5(416/590) Ro6<y6(370/590) Ro7<y7(321/590) Ro8<y8(280/590) Ro9<y9(237/590) Ro10<y10(200/590) Ro11<y11(166/590) Ro12<y12(126/590) Ro13<y13(90/590) Ro14<y14(59/590) Ro15<y15(26/590) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output y11;    //: /sn:0 {0}(360,172)(423,172)(423,175)(474,175){1}
output y13;    //: /sn:0 {0}(474,125)(395,125)(395,159)(360,159){1}
output y4;    //: /sn:0 {0}(474,378)(399,378)(399,389)(360,389){1}
output y0;    //: /sn:0 {0}(474,487)(377,487)(377,416)(360,416){1}
output y12;    //: /sn:0 {0}(360,165)(423,165)(423,149)(474,149){1}
output y8;    //: /sn:0 {0}(474,258)(375,258)(375,192)(360,192){1}
output y15;    //: /sn:0 {0}(474,79)(376,79)(376,145)(360,145){1}
output y10;    //: /sn:0 {0}(474,202)(395,202)(395,179)(360,179){1}
output y1;    //: /sn:0 {0}(474,460)(384,460)(384,409)(360,409){1}
output y2;    //: /sn:0 {0}(473,431)(392,431)(392,402)(360,402){1}
output y3;    //: /sn:0 {0}(474,404)(399,404)(399,396)(360,396){1}
output y9;    //: /sn:0 {0}(474,231)(382,231)(382,185)(360,185){1}
input [3:0] a;    //: /sn:0 {0}(#:250,503)(250,449)(250,449)(250,393){1}
//: {2}(250,392)(250,203){3}
//: {4}(250,202)(250,169){5}
//: {6}(250,168)(250,-11){7}
output y5;    //: /sn:0 {0}(474,354)(392,354)(392,382)(360,382){1}
output y7;    //: /sn:0 {0}(474,308)(377,308)(377,369)(360,369){1}
output y14;    //: /sn:0 {0}(474,101)(384,101)(384,152)(360,152){1}
output y6;    //: /sn:0 {0}(474,330)(384,330)(384,376)(360,376){1}
wire w16;    //: /sn:0 {0}(306,281)(306,430)(344,430)(344,415){1}
wire [2:0] w4;    //: /sn:0 {0}(254,169)(#:262,169)(262,169)(331,169){1}
wire [2:0] w15;    //: /sn:0 {0}(254,393)(#:262,393)(262,393)(331,393){1}
wire w5;    //: /sn:0 {0}(254,203)(279,203)(279,203)(304,203){1}
//: {2}(308,203)(344,203)(344,191){3}
//: {4}(306,205)(306,215)(306,215)(306,265){5}
//: enddecls

  assign w4 = a[2:0]; //: TAP g4 @(248,169) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  assign w15 = a[2:0]; //: TAP g3 @(248,393) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: OUT g16 (y4) @(471,378) /sn:0 /w:[ 0 ]
  //: OUT g26 (y14) @(471,101) /sn:0 /w:[ 0 ]
  //: OUT g17 (y5) @(471,354) /sn:0 /w:[ 0 ]
  //: IN g2 (a) @(250,505) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g23 (y11) @(471,175) /sn:0 /w:[ 1 ]
  _GGDECODER8 #(6, 6) g1 (.I(w15), .E(w16), .Z0(y0), .Z1(y1), .Z2(y2), .Z3(y3), .Z4(y4), .Z5(y5), .Z6(y6), .Z7(y7));   //: @(344,393) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 1 1 ] /ss:0 /do:0
  //: OUT g24 (y12) @(471,149) /sn:0 /w:[ 1 ]
  //: OUT g18 (y6) @(471,330) /sn:0 /w:[ 0 ]
  //: OUT g25 (y13) @(471,125) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g6 (.I(w5), .Z(w16));   //: @(306,271) /sn:0 /R:3 /w:[ 5 0 ]
  //: joint g7 (w5) @(306, 203) /w:[ 2 -1 1 4 ]
  //: OUT g22 (y10) @(471,202) /sn:0 /w:[ 0 ]
  //: OUT g12 (y0) @(471,487) /sn:0 /w:[ 0 ]
  assign w5 = a[3]; //: TAP g5 @(248,203) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: OUT g14 (y2) @(470,431) /sn:0 /w:[ 0 ]
  //: OUT g21 (y9) @(471,231) /sn:0 /w:[ 0 ]
  //: OUT g19 (y7) @(471,308) /sn:0 /w:[ 0 ]
  //: OUT g20 (y8) @(471,258) /sn:0 /w:[ 0 ]
  _GGDECODER8 #(6, 6) g0 (.I(w4), .E(w5), .Z0(y8), .Z1(y9), .Z2(y10), .Z3(y11), .Z4(y12), .Z5(y13), .Z6(y14), .Z7(y15));   //: @(344,169) /sn:0 /R:1 /w:[ 1 3 1 1 1 0 0 1 1 1 ] /ss:0 /do:0
  //: OUT g15 (y3) @(471,404) /sn:0 /w:[ 0 ]
  //: OUT g27 (y15) @(471,79) /sn:0 /w:[ 0 ]
  //: OUT g13 (y1) @(471,460) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU
module ALU(ALU_OUTPUT, RA, MOV, RB, LOAD, ALU_op, STR);
//: interface  /sz:(185, 240) /bd:[ Li0>RA[7:0](162/240) Li1>RB[7:0](54/240) Bi0>ALU_op[3:0](92/185) To0<LOAD(39/185) To1<MOV(94/185) To2<STR(152/185) Ro0<ALU_OUTPUT[7:0](116/240) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
reg w6;    //: /sn:0 {0}(217,317)(196,317)(196,317)(199,317){1}
output LOAD;    //: /sn:0 {0}(1045,-502)(1045,-433)(1053,-433)(1053,119)(668,119)(668,-42){1}
supply0 w50;    //: /sn:0 {0}(2206,304)(2206,289)(2172,289){1}
supply0 w39;    //: /sn:0 {0}(1351,372)(1351,346){1}
output [7:0] ALU_OUTPUT;    //: /sn:0 {0}(#:2372,395)(2384,395)(2384,557){1}
//: {2}(2386,559)(#:2410,559){3}
//: {4}(2382,559)(2295,559){5}
//: {6}(2293,557)(2293,391)(#:2258,391){7}
//: {8}(2291,559)(2084,559){9}
//: {10}(2082,557)(2082,390)(#:2063,390){11}
//: {12}(2080,559)(1905,559){13}
//: {14}(1903,557)(1903,399)(#:1891,399){15}
//: {16}(1901,559)(1686,559){17}
//: {18}(1684,557)(1684,523)(1745,523)(#:1745,381)(#:1726,381){19}
//: {20}(1682,559)(1375,559)(1375,560)(1091,560){21}
//: {22}(1089,558)(1089,431)(#:1047,431){23}
//: {24}(1087,560)(984,560){25}
//: {26}(982,558)(982,435)(#:958,435){27}
//: {28}(980,560)(901,560){29}
//: {30}(899,558)(899,443)(#:885,443){31}
//: {32}(897,560)(819,560){33}
//: {34}(817,558)(817,442)(#:798,442){35}
//: {36}(815,560)(729,560){37}
//: {38}(727,558)(727,451)(#:708,451){39}
//: {40}(725,560)(550,560){41}
//: {42}(548,558)(548,451)(#:541,451){43}
//: {44}(546,560)(426,560){45}
//: {46}(424,558)(424,450)(#:412,450){47}
//: {48}(422,560)(349,560)(349,455)(#:268,455){49}
output MOV;    //: /sn:0 {0}(1115,-479)(1115,-453)(1115,-453)(1115,-103){1}
//: {2}(1117,-101)(2364,-101)(2364,390){3}
//: {4}(1115,-99)(1115,53)(748,53)(748,-42){5}
input [7:0] RA;    //: /sn:0 {0}(#:35,262)(95,262)(95,262)(222,262){1}
//: {2}(226,262)(361,262){3}
//: {4}(365,262)(537,262){5}
//: {6}(541,262)(654,262){7}
//: {8}(#:658,262)(761,262){9}
//: {10}(#:765,262)(821,262){11}
//: {12}(#:825,262)(911,262){13}
//: {14}(#:915,262)(1000,262){15}
//: {16}(1004,262)(1038,262){17}
//: {18}(#:1042,262)(1128,262)(1128,192)(1618,192){19}
//: {20}(#:1622,192)(1787,192){21}
//: {22}(#:1791,192)(1959,192){23}
//: {24}(#:1963,192)(2130,192){25}
//: {26}(2134,192)(2341,192)(2341,395)(2356,395){27}
//: {28}(2132,194)(2132,275){29}
//: {30}(1961,194)(1961,275){31}
//: {32}(1789,194)(1789,284){33}
//: {34}(1620,194)(1620,287){35}
//: {36}(1040,264)(1040,293)(1137,293){37}
//: {38}(1002,264)(1002,306){39}
//: {40}(913,264)(913,308){41}
//: {42}(823,264)(823,300){43}
//: {44}(763,264)(763,300){45}
//: {46}(656,264)(656,302){47}
//: {48}(539,264)(#:539,269)(525,269)(525,281){49}
//: {50}(363,264)(363,303){51}
//: {52}(224,264)(224,283)(191,283)(#:191,303){53}
supply0 w44;    //: /sn:0 {0}(1412,279)(1412,316){1}
supply1 w28;    //: /sn:0 {0}(1322,220)(1322,247)(1340,247)(1340,262){1}
supply1 w35;    //: /sn:0 {0}(1368,320)(1387,320)(1387,306)(1402,306)(1402,316){1}
input [7:0] RB;    //: /sn:0 {0}(#:39,228)(190,228){1}
//: {2}(194,228)(393,228){3}
//: {4}(#:397,228)(500,228){5}
//: {6}(504,228)(686,228){7}
//: {8}(#:690,228)(766,228){9}
//: {10}(#:770,228)(826,228){11}
//: {12}(#:830,228)(995,228)(995,228)(1005,228){13}
//: {14}(1009,228)(1107,228){15}
//: {16}(#:1111,228)(1155,228)(1155,163)(1650,163){17}
//: {18}(#:1654,163)(1736,163)(1736,157)(1819,157){19}
//: {20}(#:1823,157)(1991,157){21}
//: {22}(#:1995,157)(2164,157)(2164,275){23}
//: {24}(1993,159)(1993,275){25}
//: {26}(1821,159)(1821,284){27}
//: {28}(1652,165)(1652,266)(1652,266)(1652,287){29}
//: {30}(1109,230)(1109,340)(1137,340){31}
//: {32}(1007,230)(1007,266)(1007,266)(1007,306){33}
//: {34}(828,230)(828,300){35}
//: {36}(768,230)(768,300){37}
//: {38}(688,230)(688,302){39}
//: {40}(502,230)(#:502,235)(491,235)(491,281){41}
//: {42}(395,230)(#:395,303){43}
//: {44}(192,230)(192,266)(159,266)(159,303){45}
supply1 w45;    //: /sn:0 {0}(1317,343)(1317,357)(1341,357)(1341,372){1}
reg w41;    //: /sn:0 {0}(1829,298)(1845,298)(1845,298)(1860,298){1}
supply0 w47;    //: /sn:0 {0}(2017,303)(2017,289)(2001,289){1}
input [3:0] ALU_op;    //: /sn:0 {0}(914,-377)(914,-328)(#:914,-328)(914,-233){1}
supply0 w43;    //: /sn:0 {0}(1364,234)(1364,249)(1350,249)(1350,262){1}
output STR;    //: /sn:0 {0}(1082,-493)(1082,-426)(1088,-426)(1088,90)(711,90)(711,-42){1}
reg w40;    //: /sn:0 {0}(1673,301)(1642,301)(1642,301)(1660,301){1}
wire [7:0] w13;    //: /sn:0 {0}(#:913,324)(913,435)(942,435){1}
wire [7:0] w7;    //: /sn:0 {0}(#:379,332)(379,450)(396,450){1}
wire w58;    //: /sn:0 {0}(922,-42)(922,5)(1883,5)(1883,394){1}
wire w65;    //: /sn:0 {0}(1928,276)(1928,289)(1953,289){1}
wire w34;    //: /sn:0 {0}(1287,332)(1391,332){1}
wire w59;    //: /sn:0 {0}(2055,385)(2055,-27)(889,-27)(889,-42){1}
wire w4;    //: /sn:0 {0}(103,318)(113,318)(113,303)(86,303)(86,317)(151,317){1}
wire [7:0] w25;    //: /sn:0 {0}(869,443)(825,443)(#:825,321){1}
wire w22;    //: /sn:0 {0}(498,-42)(498,14)(790,14)(790,437){1}
wire w0;    //: /sn:0 {0}(2186,386)(2186,90)(1487,90)(1487,383)(1362,383){1}
wire [7:0] w60;    //: /sn:0 {0}(2002,390)(1977,390)(#:1977,304){1}
wire w29;    //: /sn:0 {0}(578,-42)(578,-4)(950,-4)(950,430){1}
wire [7:0] w30;    //: /sn:0 {0}(#:1004,327)(1004,431)(1031,431){1}
wire w37;    //: /sn:0 {0}(1423,337)(1462,337)(1462,328){1}
wire w42;    //: /sn:0 {0}(1361,283)(1393,283)(1393,263){1}
wire [7:0] w18;    //: /sn:0 {0}(#:525,451)(491,451)(491,400){1}
wire [7:0] w19;    //: /sn:0 {0}(#:765,321)(765,442)(782,442){1}
wire [7:0] w23;    //: /sn:0 {0}(#:682,331)(682,451)(692,451){1}
wire [7:0] w54;    //: /sn:0 {0}(#:2018,390)(2025,390)(2025,390)(2047,390){1}
wire w21;    //: /sn:0 {0}(433,-42)(433,50)(533,50)(533,446){1}
wire [7:0] w24;    //: /sn:0 {0}(#:662,331)(662,369)(606,369)(606,354){1}
wire w31;    //: /sn:0 {0}(627,-42)(627,-12)(1039,-12)(1039,426){1}
wire w1;    //: /sn:0 {0}(1370,393)(1362,393){1}
wire w32;    //: /sn:0 {0}(1287,387)(1315,387)(1315,388)(1330,388){1}
wire [7:0] w53;    //: /sn:0 {0}(#:1827,399)(1834,399)(1834,399)(1875,399){1}
wire w8;    //: /sn:0 {0}(404,-42)(404,445){1}
wire [7:0] w46;    //: /sn:0 {0}(#:1636,316)(1636,381)(1710,381){1}
wire w52;    //: /sn:0 {0}(1755,276)(1755,298)(1781,298){1}
wire w27;    //: /sn:0 {0}(467,-42)(467,26)(700,26)(700,446){1}
wire w33;    //: /sn:0 {0}(1287,280)(1314,280)(1314,278)(1329,278){1}
wire [7:0] w67;    //: /sn:0 {0}(#:2194,391)(2201,391)(2201,391)(2242,391){1}
wire w14;    //: /sn:0 {0}(559,423)(525,423)(525,400){1}
wire [7:0] w49;    //: /sn:0 {0}(1811,399)(1805,399)(#:1805,313){1}
wire [7:0] w69;    //: /sn:0 {0}(2178,391)(2148,391)(#:2148,304){1}
wire [7:0] w2;    //: /sn:0 {0}(#:175,332)(175,455)(252,455){1}
wire w11;    //: /sn:0 {0}(375,-42)(375,97)(260,97)(260,450){1}
wire w48;    //: /sn:0 {0}(1592,301)(1606,301)(1606,301)(1612,301){1}
wire w74;    //: /sn:0 {0}(2106,274)(2106,289)(2124,289){1}
wire w38;    //: /sn:0 {0}(1819,394)(1819,384)(1851,384)(1851,45)(1435,45)(1435,273)(1361,273){1}
wire w61;    //: /sn:0 {0}(858,-42)(858,36)(2250,36)(2250,386){1}
wire w5;    //: /sn:0 {0}(1407,348)(1407,365)(1555,365){1}
//: {2}(1559,365)(1561,365)(1561,446)(1346,446)(1346,404){3}
//: {4}(1557,363)(1557,300)(1532,300){5}
//: {6}(1530,298)(1530,114)(782,114)(782,-42){7}
//: {8}(1528,300)(1345,300)(1345,294){9}
wire w26;    //: /sn:0 {0}(532,-42)(532,7)(877,7)(877,438){1}
wire w9;    //: /sn:0 {0}(2010,385)(2010,72)(1458,72)(1458,327)(1423,327){1}
wire w51;    //: /sn:0 {0}(822,-42)(822,-34)(1718,-34)(1718,376){1}
//: enddecls

  //: joint g8 (RA) @(539, 262) /w:[ 6 -1 5 48 ]
  //: SWITCH g4 (w6) @(235,317) /sn:0 /R:2 /w:[ 0 ] /st:0 /dn:1
  _GGBUFIF8 #(4, 6) g44 (.Z(ALU_OUTPUT), .I(w30), .E(w31));   //: @(1037,431) /sn:0 /w:[ 23 1 1 ]
  _GGBUFIF8 #(4, 6) g75 (.Z(ALU_OUTPUT), .I(w53), .E(w58));   //: @(1881,399) /sn:0 /w:[ 15 1 1 ]
  _GGBUFIF8 #(4, 6) g3 (.Z(ALU_OUTPUT), .I(w2), .E(w11));   //: @(258,455) /sn:0 /w:[ 49 1 1 ]
  //: joint g47 (RA) @(1002, 262) /w:[ 16 -1 15 38 ]
  //: joint g26 (ALU_OUTPUT) @(727, 560) /w:[ 37 38 40 -1 ]
  //: joint g90 (ALU_OUTPUT) @(2082, 559) /w:[ 9 10 12 -1 ]
  _GGBUFIF8 #(4, 6) g2 (.Z(ALU_OUTPUT), .I(w7), .E(w8));   //: @(402,450) /sn:0 /w:[ 47 1 1 ]
  _GGBUFIF8 #(4, 6) g30 (.Z(ALU_OUTPUT), .I(w19), .E(w22));   //: @(788,442) /sn:0 /w:[ 35 1 1 ]
  _GGBUFIF8 #(4, 6) g74 (.Z(w53), .I(w49), .E(w38));   //: @(1817,399) /sn:0 /w:[ 0 0 0 ]
  //: joint g91 (ALU_OUTPUT) @(2293, 559) /w:[ 5 6 8 -1 ]
  //: OUT g92 (ALU_OUTPUT) @(2407,559) /sn:0 /w:[ 3 ]
  _GGMUL8 #(124) g1 (.A(RA), .B(RB), .P(w7));   //: @(379,319) /sn:0 /w:[ 51 43 0 ]
  //: joint g24 (ALU_OUTPUT) @(548, 560) /w:[ 41 42 44 -1 ]
  _GGBUFIF8 #(4, 6) g39 (.Z(ALU_OUTPUT), .I(w13), .E(w29));   //: @(948,435) /sn:0 /w:[ 27 1 1 ]
  _GGBUFIF8 #(4, 6) g77 (.Z(w54), .I(w60), .E(w9));   //: @(2008,390) /sn:0 /w:[ 0 0 0 ]
  //: joint g86 (RA) @(1961, 192) /w:[ 24 -1 23 30 ]
  //: joint g29 (RB) @(688, 228) /w:[ 8 -1 7 38 ]
  //: VDD g60 (w45) @(1328,343) /sn:0 /w:[ 0 ]
  //: IN g51 (RA) @(33,262) /sn:0 /w:[ 0 ]
  _GGBUFIF8 #(4, 6) g18 (.Z(ALU_OUTPUT), .I(w18), .E(w21));   //: @(531,451) /sn:0 /w:[ 43 0 1 ]
  //: joint g70 (RB) @(1109, 228) /w:[ 16 -1 15 30 ]
  //: joint g82 (RA) @(1620, 192) /w:[ 20 -1 19 34 ]
  //: LED g10 (w14) @(566,423) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: joint g25 (ALU_OUTPUT) @(424, 560) /w:[ 45 46 48 -1 ]
  //: joint g65 (w5) @(1557, 365) /w:[ 2 4 1 -1 ]
  //: LED g94 (w52) @(1755,269) /sn:0 /w:[ 0 ] /type:0
  //: LED g64 (w1) @(1377,393) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: joint g49 (RA) @(224, 262) /w:[ 2 -1 1 52 ]
  //: LED g72 (w48) @(1585,301) /sn:0 /R:1 /w:[ 0 ] /type:0
  final_sub g6 (.A(RA), .B(RB), .COUT(w14), .S(w18));   //: @(457, 282) /sz:(103, 117) /R:3 /sn:0 /p:[ Ti0>49 Ti1>41 Bo0<1 Bo1<1 ]
  //: joint g50 (RB) @(192, 228) /w:[ 2 -1 1 44 ]
  //: joint g9 (RB) @(502, 228) /w:[ 6 -1 5 40 ]
  //: joint g7 (RA) @(363, 262) /w:[ 4 -1 3 50 ]
  _GGBUFIF8 #(4, 6) g35 (.Z(ALU_OUTPUT), .I(w25), .E(w26));   //: @(875,443) /sn:0 /w:[ 31 0 1 ]
  //: GROUND g56 (w43) @(1364,228) /sn:0 /R:2 /w:[ 0 ]
  //: GROUND g58 (w39) @(1351,340) /sn:0 /R:2 /w:[ 1 ]
  _GGBUFIF8 #(4, 6) g68 (.Z(ALU_OUTPUT), .I(w46), .E(w51));   //: @(1716,381) /sn:0 /w:[ 19 1 1 ]
  _GGADD8 #(68, 70, 62, 64) g73 (.A(RA), .B(RB), .S(w49), .CI(w41), .CO(w52));   //: @(1805,300) /sn:0 /w:[ 33 27 1 0 1 ]
  //: joint g31 (ALU_OUTPUT) @(817, 560) /w:[ 33 34 36 -1 ]
  //: VDD g59 (w28) @(1333,220) /sn:0 /w:[ 0 ]
  //: SWITCH g71 (w40) @(1691,301) /sn:0 /R:2 /w:[ 0 ] /st:0 /dn:1
  //: LED g98 (w74) @(2106,267) /sn:0 /w:[ 0 ] /type:0
  //: OUT g102 (MOV) @(1115,-476) /sn:0 /R:1 /w:[ 0 ]
  _GGADD8 #(68, 70, 62, 64) g67 (.A(RA), .B(RB), .S(w46), .CI(w40), .CO(w48));   //: @(1636,303) /sn:0 /w:[ 35 29 0 1 1 ]
  //: joint g85 (RB) @(1821, 157) /w:[ 20 -1 19 26 ]
  //: joint g87 (RB) @(1993, 157) /w:[ 22 -1 21 24 ]
  //: joint g83 (RB) @(1652, 163) /w:[ 18 -1 17 28 ]
  //: GROUND g99 (w50) @(2206,310) /sn:0 /w:[ 0 ]
  //: joint g33 (RA) @(763, 262) /w:[ 10 -1 9 44 ]
  //: joint g36 (ALU_OUTPUT) @(899, 560) /w:[ 29 30 32 -1 ]
  _GGXOR2x8 #(8) g41 (.I0(RB), .I1(RA), .Z(w30));   //: @(1004,317) /sn:0 /R:3 /w:[ 33 39 0 ]
  //: joint g45 (ALU_OUTPUT) @(1089, 560) /w:[ 21 22 24 -1 ]
  _GGFF #(10, 10, 20) g54 (.Q(w9), ._Q(w37), .D(w34), .EN(w44), .CLR(w35), .CK(w5));   //: @(1407,332) /sn:0 /w:[ 1 0 1 1 1 0 ] /mi:0
  //: joint g40 (ALU_OUTPUT) @(982, 560) /w:[ 25 26 28 -1 ]
  //: joint g42 (RA) @(913, 262) /w:[ 14 -1 13 40 ]
  //: IN g52 (RB) @(37,228) /sn:0 /w:[ 0 ]
  //: joint g69 (RA) @(1040, 262) /w:[ 18 -1 17 36 ]
  _GGADD8 #(68, 70, 62, 64) g81 (.A(RA), .B(RB), .S(w69), .CI(w50), .CO(w74));   //: @(2148,291) /sn:0 /w:[ 29 23 1 1 1 ]
  //: joint g66 (w5) @(1530, 300) /w:[ 5 6 8 -1 ]
  //: joint g12 (RB) @(395, 228) /w:[ 4 -1 3 42 ]
  //: joint g28 (RA) @(656, 262) /w:[ 8 -1 7 46 ]
  //: joint g34 (RB) @(768, 228) /w:[ 10 -1 9 36 ]
  comp g46 (.a(RA), .b(RB), .et(w34), .gt(w33), .lt(w32));   //: @(1138, 246) /sz:(148, 189) /sn:0 /p:[ Li0>37 Li1>31 Ro0<0 Ro1<0 Ro2<0 ]
  //: GROUND g57 (w44) @(1412,273) /sn:0 /R:2 /w:[ 0 ]
  //: joint g14 (ALU_OUTPUT) @(2384, 559) /w:[ 2 1 4 -1 ]
  //: joint g11 (RA) @(2132, 192) /w:[ 26 -1 25 28 ]
  //: LED g5 (w4) @(96,318) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: joint g84 (RA) @(1789, 192) /w:[ 22 -1 21 32 ]
  //: LED g96 (w65) @(1928,269) /sn:0 /w:[ 0 ] /type:0
  _GGDIV8 #(236, 236) g19 (.A(RA), .B(RB), .Q(w23), .R(w24));   //: @(672,318) /sn:0 /w:[ 47 39 0 0 ]
  _GGBUFIF8 #(4, 6) g21 (.Z(ALU_OUTPUT), .I(w23), .E(w27));   //: @(698,451) /sn:0 /w:[ 39 1 1 ]
  //: VDD g61 (w35) @(1368,309) /sn:0 /R:1 /w:[ 0 ]
  //: LED g20 (w24) @(606,347) /sn:0 /w:[ 1 ] /type:1
  _GGOR2x8 #(6) g32 (.I0(RB), .I1(RA), .Z(w25));   //: @(825,311) /sn:0 /R:3 /w:[ 35 43 1 ]
  _GGADD8 #(68, 70, 62, 64) g78 (.A(RA), .B(RB), .S(w60), .CI(w47), .CO(w65));   //: @(1977,291) /sn:0 /w:[ 31 25 1 1 1 ]
  _GGBUFIF8 #(4, 6) g79 (.Z(ALU_OUTPUT), .I(w67), .E(w61));   //: @(2248,391) /sn:0 /w:[ 7 1 1 ]
  //: LED g63 (w37) @(1462,321) /sn:0 /w:[ 1 ] /type:0
  //: GROUND g97 (w47) @(2017,309) /sn:0 /w:[ 0 ]
  //: OUT g100 (LOAD) @(1045,-499) /sn:0 /R:1 /w:[ 0 ]
  //: IN g93 (ALU_op) @(914,-379) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (MOV) @(1115, -101) /w:[ 2 1 -1 4 ]
  _GGADD8 #(68, 70, 62, 64) g0 (.A(RB), .B(RA), .S(w2), .CI(w6), .CO(w4));   //: @(175,319) /sn:0 /w:[ 45 53 0 1 1 ]
  //: joint g38 (RA) @(823, 262) /w:[ 12 -1 11 42 ]
  //: joint g43 (RB) @(828, 228) /w:[ 12 -1 11 34 ]
  //: joint g89 (ALU_OUTPUT) @(1903, 559) /w:[ 13 14 16 -1 ]
  //: OUT g101 (STR) @(1082,-490) /sn:0 /R:1 /w:[ 0 ]
  _GGAND2x8 #(6) g27 (.I0(RB), .I1(RA), .Z(w19));   //: @(765,311) /sn:0 /R:3 /w:[ 37 45 0 ]
  //: joint g48 (RB) @(1007, 228) /w:[ 14 -1 13 32 ]
  _GGNBUF8 #(2) g37 (.I(RA), .Z(w13));   //: @(913,314) /sn:0 /R:3 /w:[ 41 0 ]
  //: LED g62 (w42) @(1393,256) /sn:0 /w:[ 1 ] /type:0
  _GGFF #(10, 10, 20) g55 (.Q(w38), ._Q(w42), .D(w33), .EN(w43), .CLR(w28), .CK(w5));   //: @(1345,278) /sn:0 /w:[ 1 0 1 1 1 9 ] /mi:0
  _GGBUFIF8 #(4, 6) g80 (.Z(w67), .I(w69), .E(w0));   //: @(2184,391) /sn:0 /w:[ 0 0 0 ]
  //: joint g88 (ALU_OUTPUT) @(1684, 559) /w:[ 17 18 20 -1 ]
  //: SWITCH g95 (w41) @(1878,298) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  dec_4to16 DECODER (.a(ALU_op), .y0(w11), .y1(w8), .y2(w21), .y3(w27), .y4(w22), .y5(w26), .y6(w29), .y7(w31), .y8(LOAD), .y9(STR), .y10(MOV), .y11(w5), .y12(w51), .y13(w61), .y14(w59), .y15(w58));   //: @(358, -232) /sz:(590, 189) /R:3 /p:[ Ti0>1 Bo0<0 Bo1<0 Bo2<0 Bo3<0 Bo4<0 Bo5<0 Bo6<0 Bo7<0 Bo8<1 Bo9<1 Bo10<5 Bo11<7 Bo12<0 Bo13<0 Bo14<1 Bo15<0 ]
  _GGBUFIF8 #(4, 6) g13 (.Z(ALU_OUTPUT), .I(RA), .E(MOV));   //: @(2362,395) /sn:0 /w:[ 0 27 3 ]
  _GGFF #(10, 10, 20) g53 (.Q(w0), ._Q(w1), .D(w32), .EN(w39), .CLR(w45), .CK(w5));   //: @(1346,388) /sn:0 /w:[ 1 1 1 0 1 3 ] /mi:0
  _GGBUFIF8 #(4, 6) g76 (.Z(ALU_OUTPUT), .I(w54), .E(w59));   //: @(2053,390) /sn:0 /w:[ 11 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin F_Add
module F_Add(cout, b, sum, cin, a);
//: interface  /sz:(93, 64) /bd:[ Li0>cin(48/64) Li1>b(32/64) Li2>a(16/64) Ro0<sum(32/64) Ro1<cout(16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(140,144)(149,144)(149,144)(157,144){1}
//: {2}(161,144)(171,144)(171,144)(179,144){3}
//: {4}(159,146)(159,285)(262,285){5}
input cin;    //: /sn:0 {0}(132,204)(238,204)(238,204)(208,204){1}
//: {2}(212,204)(248,204)(248,147)(261,147){3}
//: {4}(210,206)(210,230)(261,230){5}
output sum;    //: /sn:0 {0}(282,145)(378,145)(378,145)(393,145){1}
output cout;    //: /sn:0 {0}(378,256)(372,256)(372,256)(392,256){1}
input a;    //: /sn:0 {0}(125,139)(138,139)(138,139)(146,139){1}
//: {2}(150,139)(179,139){3}
//: {4}(148,141)(148,290)(262,290){5}
wire w0;    //: /sn:0 {0}(200,142)(219,142){1}
//: {2}(223,142)(248,142)(248,142)(261,142){3}
//: {4}(221,144)(221,225)(261,225){5}
wire w2;    //: /sn:0 {0}(282,228)(342,228)(342,253)(357,253){1}
wire w5;    //: /sn:0 {0}(283,288)(342,288)(342,258)(357,258){1}
//: enddecls

  //: OUT g8 (cout) @(389,256) /sn:0 /w:[ 1 ]
  _GGXOR2 #(8) g4 (.I0(a), .I1(b), .Z(w0));   //: @(190,142) /sn:0 /w:[ 3 3 0 ]
  _GGXOR2 #(8) g3 (.I0(w0), .I1(cin), .Z(sum));   //: @(272,145) /sn:0 /w:[ 3 3 0 ]
  _GGOR2 #(6) g2 (.I0(w2), .I1(w5), .Z(cout));   //: @(368,256) /sn:0 /w:[ 1 1 0 ]
  _GGAND2 #(6) g1 (.I0(b), .I1(a), .Z(w5));   //: @(273,288) /sn:0 /w:[ 5 5 0 ]
  //: joint g10 (w0) @(221, 142) /w:[ 2 -1 1 4 ]
  //: IN g6 (b) @(138,144) /sn:0 /w:[ 0 ]
  //: OUT g9 (sum) @(390,145) /sn:0 /w:[ 1 ]
  //: IN g7 (cin) @(130,204) /sn:0 /w:[ 0 ]
  //: joint g12 (b) @(159, 144) /w:[ 2 -1 1 4 ]
  //: joint g11 (cin) @(210, 204) /w:[ 2 -1 1 4 ]
  //: IN g5 (a) @(123,139) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g0 (.I0(w0), .I1(cin), .Z(w2));   //: @(272,228) /sn:0 /w:[ 5 5 0 ]
  //: joint g13 (a) @(148, 139) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin demux
module demux(D1, D0, RF, RY, PC);
//: interface  /sz:(112, 102) /bd:[ Ti0>D1(63/112) Ti1>D0(35/112) Ri0>RY[7:0](16/102) Lo0<RF[7:0](70/102) Lo1<PC[7:0](25/102) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] PC;    //: /sn:0 {0}(#:226,375)(230,375)(230,155)(141,155)(141,195)(87,195){1}
input D1;    //: /sn:0 {0}(365,-10)(365,21)(355,21)(355,309){1}
//: {2}(357,311)(413,311)(413,296)(428,296){3}
//: {4}(355,313)(355,371){5}
input [7:0] RY;    //: /sn:0 {0}(#:490,5)(490,66)(673,66)(673,464)(130,464)(130,338)(175,338){1}
//: {2}(179,338)(327,338){3}
//: {4}(331,338)(462,338)(462,374)(#:475,374){5}
//: {6}(#:329,340)(329,376)(347,376){7}
//: {8}(177,340)(177,375)(#:210,375){9}
input D0;    //: /sn:0 {0}(252,-1)(280,-1)(280,41)(218,41)(218,278){1}
//: {2}(220,280)(413,280)(413,291)(428,291){3}
//: {4}(218,282)(218,370){5}
output [7:0] RF;    //: /sn:0 {0}(105,247)(408,247)(408,376)(#:363,376){1}
wire w94;    //: /sn:0 {0}(449,294)(483,294)(483,369){1}
wire [7:0] w92;    //: /sn:0 {0}(525,174)(525,374)(#:491,374){1}
//: enddecls

  //: IN g4 (D1) @(365,-12) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (D0) @(250,-1) /sn:0 /w:[ 0 ]
  //: LED g2 (w92) @(525,167) /sn:0 /w:[ 0 ] /type:1
  //: OUT g1 (RF) @(108,247) /sn:0 /R:2 /w:[ 0 ]
  //: joint g220 (D1) @(355, 311) /w:[ 2 1 -1 4 ]
  _GGBUFIF8 #(4, 6) g216 (.Z(RF), .I(RY), .E(D1));   //: @(353,376) /sn:0 /w:[ 1 7 5 ]
  _GGBUFIF8 #(4, 6) g217 (.Z(w92), .I(RY), .E(w94));   //: @(481,374) /sn:0 /w:[ 1 5 1 ]
  //: IN g5 (RY) @(490,3) /sn:0 /R:3 /w:[ 0 ]
  _GGNOR2 #(4) g221 (.I0(D0), .I1(D1), .Z(w94));   //: @(439,294) /sn:0 /w:[ 3 3 0 ]
  //: joint g219 (RY) @(329, 338) /w:[ 4 -1 3 6 ]
  //: OUT g0 (PC) @(90,195) /sn:0 /R:2 /w:[ 1 ]
  _GGBUFIF8 #(4, 6) g215 (.Z(PC), .I(RY), .E(D0));   //: @(216,375) /sn:0 /w:[ 0 9 5 ]
  //: joint g147 (RY) @(177, 338) /w:[ 2 -1 1 8 ]
  //: joint g218 (D0) @(218, 280) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin register_file
module register_file(ra_s, A, C, CLK, Add_A, rc_s, Add_B, B, Add_C, CLR, rb_s);
//: interface  /sz:(155, 434) /bd:[ Ti0>C[7:0](80/155) Li0>Add_A[2:0](74/434) Li1>Add_B[2:0](118/434) Li2>ra_s(190/434) Li3>rb_s(223/434) Li4>rc_s(252/434) Li5>CLK(311/434) Li6>CLR(361/434) Ri0>Add_C[2:0](137/434) Bo0<A[7:0](20/155) Bo1<B[7:0](134/155) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] B;    //: /sn:0 {0}(#:865,379)(652,379){1}
//: {2}(650,377)(650,311){3}
//: {4}(650,307)(650,208){5}
//: {6}(650,204)(650,94){7}
//: {8}(650,90)(650,-8)(#:545,-8){9}
//: {10}(648,92)(603,92)(603,92)(#:556,92){11}
//: {12}(648,206)(602,206)(602,206)(#:556,206){13}
//: {14}(648,309)(604,309)(604,309)(#:556,309){15}
//: {16}(650,381)(650,398){17}
//: {18}(648,400)(#:556,400){19}
//: {20}(650,402)(650,447)(650,447)(650,491){21}
//: {22}(648,493)(601,493)(601,493)(#:556,493){23}
//: {24}(650,495)(650,600){25}
//: {26}(648,602)(597,602)(597,602)(#:556,602){27}
//: {28}(650,604)(650,725)(#:562,725){29}
supply0 w4;    //: /sn:0 {0}(498,686)(498,667){1}
//: {2}(498,663)(498,564){3}
//: {4}(498,560)(498,509)(498,509)(498,458){5}
//: {6}(498,454)(498,361){7}
//: {8}(498,357)(498,261){9}
//: {10}(498,257)(498,166){11}
//: {12}(498,162)(498,56){13}
//: {14}(498,52)(498,-48)(460,-48){15}
//: {16}(496,54)(466,54){17}
//: {18}(496,164)(462,164){19}
//: {20}(496,259)(466,259){21}
//: {22}(496,359)(481,359)(481,359)(466,359){23}
//: {24}(496,456)(466,456){25}
//: {26}(496,562)(468,562){27}
//: {28}(496,665)(469,665){29}
output [7:0] A;    //: /sn:0 {0}(#:868,279)(707,279){1}
//: {2}(705,277)(705,265){3}
//: {4}(705,261)(705,211)(705,211)(705,161){5}
//: {6}(705,157)(705,47){7}
//: {8}(705,43)(705,-59)(#:535,-59){9}
//: {10}(703,45)(#:556,45){11}
//: {12}(703,159)(#:553,159){13}
//: {14}(703,263)(693,263)(693,263)(#:556,263){15}
//: {16}(705,281)(705,358){17}
//: {18}(703,360)(#:556,360){19}
//: {20}(705,362)(705,451){21}
//: {22}(703,453)(#:556,453){23}
//: {24}(705,455)(705,502)(705,502)(705,549){25}
//: {26}(703,551)(#:557,551){27}
//: {28}(705,553)(705,685)(#:562,685){29}
input ra_s;    //: /sn:0 {0}(508,-368)(508,-258)(543,-258){1}
input rb_s;    //: /sn:0 {0}(602,-328)(602,-281)(627,-281)(627,-208)(649,-208){1}
input [2:0] Add_B;    //: /sn:0 {0}(#:673,-315)(673,-221){1}
input [2:0] Add_A;    //: /sn:0 {0}(#:567,-358)(567,-271){1}
input rc_s;    //: /sn:0 {0}(10,-204)(29,-204)(29,-217)(44,-217)(44,-259)(72,-259){1}
input CLR;    //: /sn:0 {0}(460,-58)(483,-58){1}
//: {2}(485,-60)(485,-193)(399,-193)(399,-239)(440,-239)(440,-217)(458,-217){3}
//: {4}(485,-56)(485,42){5}
//: {6}(483,44)(466,44){7}
//: {8}(485,46)(485,152){9}
//: {10}(483,154)(462,154){11}
//: {12}(485,156)(485,247){13}
//: {14}(483,249)(466,249){15}
//: {16}(485,251)(485,347){17}
//: {18}(483,349)(475,349)(475,349)(466,349){19}
//: {20}(485,351)(485,444){21}
//: {22}(483,446)(466,446){23}
//: {24}(485,448)(485,499)(485,499)(485,550){25}
//: {26}(483,552)(468,552){27}
//: {28}(485,554)(485,655)(469,655){29}
input [7:0] C;    //: /sn:0 {0}(430,650)(430,645)(#:320,645){1}
//: {2}(318,643)(318,531){3}
//: {4}(#:320,529)(429,529)(429,547){5}
//: {6}(318,527)(318,481)(318,481)(318,435){7}
//: {8}(#:320,433)(427,433)(427,441){9}
//: {10}(318,431)(318,334){11}
//: {12}(#:320,332)(427,332)(427,344){13}
//: {14}(318,330)(318,235){15}
//: {16}(#:320,233)(427,233)(427,244){17}
//: {18}(318,231)(318,139){19}
//: {20}(#:320,137)(423,137)(423,149){21}
//: {22}(318,135)(318,26){23}
//: {24}(320,24)(427,24)(427,39){25}
//: {26}(318,22)(318,-113)(421,-113)(421,-63){27}
//: {28}(318,647)(318,781)(#:909,781){29}
input CLK;    //: /sn:0 {0}(179,-311)(265,-311)(265,-286)(232,-286)(232,-205)(134,-205)(134,-53){1}
//: {2}(136,-51)(148,-51){3}
//: {4}(134,-49)(134,49){5}
//: {6}(136,51)(147,51){7}
//: {8}(134,53)(134,159){9}
//: {10}(136,161)(147,161){11}
//: {12}(134,163)(134,254){13}
//: {14}(136,256)(147,256){15}
//: {16}(134,258)(134,354){17}
//: {18}(136,356)(147,356){19}
//: {20}(134,358)(134,451){21}
//: {22}(136,453)(147,453){23}
//: {24}(134,455)(134,506)(134,506)(134,557){25}
//: {26}(136,559)(147,559){27}
//: {28}(134,561)(134,662)(147,662){29}
input [2:0] Add_C;    //: /sn:0 {0}(#:96,-335)(96,-272){1}
wire [7:0] w16;    //: /sn:0 {0}(#:427,365)(427,381)(427,381)(427,398){1}
//: {2}(429,400)(517,400){3}
//: {4}(521,400)(540,400){5}
//: {6}(#:519,398)(519,360)(540,360){7}
//: {8}(#:425,400)(357,400)(357,378){9}
wire [7:0] w6;    //: /sn:0 {0}(#:540,206)(530,206){1}
//: {2}(#:528,204)(528,159)(537,159){3}
//: {4}(526,206)(425,206){5}
//: {6}(423,204)(#:423,170){7}
//: {8}(#:421,206)(357,206)(357,184){9}
wire w58;    //: /sn:0 {0}(656,-192)(656,124)(563,124)(563,77)(548,77)(548,87){1}
wire w65;    //: /sn:0 {0}(590,-242)(590,708)(565,708)(565,673)(554,673)(554,680){1}
wire w34;    //: /sn:0 {0}(557,-242)(557,144)(545,144)(545,154){1}
wire w88;    //: /sn:0 {0}(80,-243)(80,46)(147,46){1}
wire w59;    //: /sn:0 {0}(583,-242)(583,534)(549,534)(549,546){1}
wire w25;    //: /sn:0 {0}(168,451)(218,451)(218,451)(390,451){1}
wire w39;    //: /sn:0 {0}(563,-242)(563,246)(548,246)(548,258){1}
wire [7:0] w72;    //: /sn:0 {0}(#:429,568)(429,600){1}
//: {2}(431,602)(517,602){3}
//: {4}(521,602)(540,602){5}
//: {6}(#:519,600)(519,551)(541,551){7}
//: {8}(#:427,602)(357,602)(357,585){9}
wire w101;    //: /sn:0 {0}(86,-243)(86,156)(147,156){1}
wire [7:0] w36;    //: /sn:0 {0}(#:430,671)(430,723){1}
//: {2}(432,725)(533,725){3}
//: {4}(537,725)(546,725){5}
//: {6}(#:535,723)(535,685)(546,685){7}
//: {8}(#:428,725)(357,725)(357,690){9}
wire w20;    //: /sn:0 {0}(168,354)(390,354){1}
wire w30;    //: /sn:0 {0}(168,557)(227,557)(227,557)(392,557){1}
wire w73;    //: /sn:0 {0}(689,-192)(689,637)(563,637)(563,587)(548,587)(548,597){1}
wire [7:0] w63;    //: /sn:0 {0}(#:427,265)(427,307){1}
//: {2}(429,309)(521,309){3}
//: {4}(525,309)(540,309){5}
//: {6}(#:523,307)(523,263)(540,263){7}
//: {8}(#:425,309)(357,309)(357,283){9}
wire w10;    //: /sn:0 {0}(168,159)(238,159)(238,159)(386,159){1}
wire [7:0] w23;    //: /sn:0 {0}(#:421,-42)(421,-10){1}
//: {2}(423,-8)(522,-8){3}
//: {4}(526,-8)(529,-8){5}
//: {6}(524,-10)(524,-30)(509,-30)(509,-59)(519,-59){7}
//: {8}(#:419,-8)(373,-8)(373,-22){9}
wire w70;    //: /sn:0 {0}(683,-192)(683,528)(563,528)(563,478)(548,478)(548,488){1}
wire w91;    //: /sn:0 {0}(100,-243)(100,351)(147,351){1}
wire [7:0] w21;    //: /sn:0 {0}(#:427,462)(427,477)(427,477)(427,491){1}
//: {2}(429,493)(520,493){3}
//: {4}(524,493)(540,493){5}
//: {6}(#:522,491)(522,453)(540,453){7}
//: {8}(#:425,493)(357,493)(357,474){9}
wire [7:0] w1;    //: /sn:0 {0}(#:540,92)(530,92){1}
//: {2}(#:528,90)(528,45)(540,45){3}
//: {4}(526,92)(451,92)(451,92)(429,92){5}
//: {6}(427,90)(#:427,60){7}
//: {8}(#:425,92)(357,92)(357,78){9}
wire w31;    //: /sn:0 {0}(548,40)(548,26)(550,26)(550,-242){1}
wire w104;    //: /sn:0 {0}(93,-243)(93,251)(147,251){1}
wire w116;    //: /sn:0 {0}(120,-243)(120,657)(147,657){1}
wire w53;    //: /sn:0 {0}(577,-242)(577,435)(548,435)(548,448){1}
wire w110;    //: /sn:0 {0}(106,-243)(106,448)(147,448){1}
wire w46;    //: /sn:0 {0}(570,-242)(570,347)(548,347)(548,355){1}
wire w95;    //: /sn:0 {0}(73,-243)(73,-56)(148,-56){1}
wire w27;    //: /sn:0 {0}(527,-64)(527,-80)(543,-80)(543,-242){1}
wire w67;    //: /sn:0 {0}(676,-192)(676,434)(563,434)(563,385)(548,385)(548,395){1}
wire w113;    //: /sn:0 {0}(113,-243)(113,554)(147,554){1}
wire w35;    //: /sn:0 {0}(169,-53)(384,-53){1}
wire w15;    //: /sn:0 {0}(168,254)(226,254)(226,254)(390,254){1}
wire w5;    //: /sn:0 {0}(168,49)(233,49)(233,49)(390,49){1}
wire w55;    //: /sn:0 {0}(649,-192)(649,24)(552,24)(552,-23)(537,-23)(537,-13){1}
wire w61;    //: /sn:0 {0}(663,-192)(663,238)(563,238)(563,191)(548,191)(548,201){1}
wire w64;    //: /sn:0 {0}(669,-192)(669,343)(563,343)(563,294)(548,294)(548,304){1}
wire w76;    //: /sn:0 {0}(696,-192)(696,760)(569,760)(569,710)(554,710)(554,720){1}
wire w40;    //: /sn:0 {0}(168,660)(221,660)(221,660)(393,660){1}
//: enddecls

  //: joint g44 (B) @(650, 206) /w:[ -1 6 12 5 ]
  //: joint g75 (w63) @(427, 309) /w:[ 2 1 8 -1 ]
  _GGAND2 #(6) g178 (.I0(w110), .I1(CLK), .Z(w25));   //: @(158,451) /sn:0 /w:[ 1 23 0 ]
  _GGREG8 #(10, 10, 20) g8 (.Q(w36), .D(C), .EN(w4), .CLR(~CLR), .CK(w40));   //: @(430,660) /sn:0 /w:[ 0 0 29 29 1 ]
  _GGREG8 #(10, 10, 20) g4 (.Q(w16), .D(C), .EN(w4), .CLR(~CLR), .CK(w20));   //: @(427,354) /sn:0 /w:[ 0 13 23 19 1 ]
  _GGBUFIF8 #(4, 6) g16 (.Z(B), .I(w16), .E(w67));   //: @(546,400) /sn:0 /w:[ 19 5 1 ]
  _GGREG8 #(10, 10, 20) g3 (.Q(w63), .D(C), .EN(w4), .CLR(~CLR), .CK(w15));   //: @(427,254) /sn:0 /w:[ 0 17 21 15 1 ]
  //: joint g47 (B) @(650, 400) /w:[ -1 17 18 20 ]
  //: joint g182 (CLK) @(134, -51) /w:[ 2 1 -1 4 ]
  //: joint g26 (C) @(318, 529) /w:[ 4 6 -1 3 ]
  _GGBUFIF8 #(4, 6) g90 (.Z(A), .I(w6), .E(w34));   //: @(543,159) /sn:0 /w:[ 13 3 1 ]
  //: joint g109 (A) @(705, 551) /w:[ -1 25 26 28 ]
  _GGBUFIF8 #(4, 6) g17 (.Z(B), .I(w21), .E(w70));   //: @(546,493) /sn:0 /w:[ 23 5 1 ]
  _GGREG8 #(10, 10, 20) g2 (.Q(w6), .D(C), .EN(w4), .CLR(~CLR), .CK(w10));   //: @(423,159) /sn:0 /w:[ 7 21 19 11 1 ]
  _GGAND2 #(6) g174 (.I0(w88), .I1(CLK), .Z(w5));   //: @(158,49) /sn:0 /w:[ 1 7 0 ]
  //: joint g23 (C) @(318, 233) /w:[ 16 18 -1 15 ]
  _GGBUFIF8 #(4, 6) g91 (.Z(A), .I(w63), .E(w39));   //: @(546,263) /sn:0 /w:[ 15 7 1 ]
  //: joint g30 (CLR) @(485, 154) /w:[ -1 9 10 12 ]
  //: joint g74 (w6) @(423, 206) /w:[ 5 6 8 -1 ]
  _GGBUFIF8 #(4, 6) g92 (.Z(A), .I(w16), .E(w46));   //: @(546,360) /sn:0 /w:[ 19 7 1 ]
  //: joint g24 (C) @(318, 332) /w:[ 12 14 -1 11 ]
  //: joint g39 (w4) @(498, 456) /w:[ -1 6 24 5 ]
  //: joint g104 (A) @(705, 45) /w:[ -1 8 10 7 ]
  _GGREG8 #(10, 10, 20) g1 (.Q(w1), .D(C), .EN(w4), .CLR(~CLR), .CK(w5));   //: @(427,49) /sn:0 /w:[ 7 25 17 7 1 ]
  //: joint g77 (w21) @(427, 493) /w:[ 2 1 8 -1 ]
  //: joint g183 (CLK) @(134, 51) /w:[ 6 5 -1 8 ]
  //: joint g29 (CLR) @(485, 44) /w:[ -1 5 6 8 ]
  _GGDECODER8 #(6, 6) g168 (.I(Add_B), .E(rb_s), .Z0(w55), .Z1(w58), .Z2(w61), .Z3(w64), .Z4(w67), .Z5(w70), .Z6(w73), .Z7(w76));   //: @(673,-208) /sn:0 /w:[ 1 1 0 0 0 0 0 0 0 0 ] /ss:0 /do:0
  _GGAND2 #(6) g179 (.I0(w113), .I1(CLK), .Z(w30));   //: @(158,557) /sn:0 /w:[ 1 27 0 ]
  //: IN g51 (ra_s) @(508,-370) /sn:0 /R:3 /w:[ 0 ]
  _GGBUFIF8 #(4, 6) g18 (.Z(B), .I(w72), .E(w73));   //: @(546,602) /sn:0 /w:[ 27 5 1 ]
  //: LED g70 (w72) @(357,578) /sn:0 /w:[ 9 ] /type:1
  _GGBUFIF8 #(4, 6) g94 (.Z(A), .I(w72), .E(w59));   //: @(547,551) /sn:0 /w:[ 27 7 1 ]
  //: joint g25 (C) @(318, 433) /w:[ 8 10 -1 7 ]
  //: LED g65 (w1) @(357,71) /sn:0 /w:[ 9 ] /type:1
  //: joint g103 (w36) @(535, 725) /w:[ 4 6 3 -1 ]
  //: OUT g10 (A) @(865,279) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g173 (.I0(w95), .I1(CLK), .Z(w35));   //: @(159,-53) /sn:0 /w:[ 1 3 0 ]
  //: joint g107 (A) @(705, 360) /w:[ -1 17 18 20 ]
  //: LED g64 (w23) @(373,-29) /sn:0 /w:[ 9 ] /type:1
  //: joint g188 (CLK) @(134, 559) /w:[ 26 25 -1 28 ]
  //: joint g184 (CLK) @(134, 161) /w:[ 10 9 -1 12 ]
  _GGDECODER8 #(6, 6) g172 (.I(Add_C), .E(rc_s), .Z0(w95), .Z1(w88), .Z2(w101), .Z3(w104), .Z4(w91), .Z5(w110), .Z6(w113), .Z7(w116));   //: @(96,-259) /sn:0 /w:[ 1 1 0 0 0 0 0 0 0 0 ] /ss:0 /do:0
  //: joint g49 (B) @(650, 602) /w:[ -1 25 26 28 ]
  //: joint g72 (w36) @(430, 725) /w:[ 2 1 8 -1 ]
  //: joint g185 (CLK) @(134, 256) /w:[ 14 13 -1 16 ]
  _GGREG8 #(10, 10, 20) g6 (.Q(w72), .D(C), .EN(w4), .CLR(~CLR), .CK(w30));   //: @(429,557) /sn:0 /w:[ 0 5 27 27 1 ]
  //: IN g50 (C) @(911,781) /sn:0 /R:2 /w:[ 29 ]
  //: joint g73 (w1) @(427, 92) /w:[ 5 6 8 -1 ]
  //: LED g68 (w16) @(357,371) /sn:0 /w:[ 9 ] /type:1
  _GGREG8 #(10, 10, 20) g7 (.Q(w23), .D(C), .EN(w4), .CLR(~CLR), .CK(w35));   //: @(421,-53) /sn:0 /w:[ 0 27 15 0 1 ]
  //: GROUND g35 (w4) @(498,692) /sn:0 /w:[ 0 ]
  //: joint g9 (B) @(650, 379) /w:[ 1 2 -1 16 ]
  //: IN g56 (CLK) @(177,-311) /sn:0 /w:[ 0 ]
  //: joint g186 (CLK) @(134, 356) /w:[ 18 17 -1 20 ]
  //: joint g102 (w72) @(519, 602) /w:[ 4 6 3 -1 ]
  //: LED g71 (w36) @(357,683) /sn:0 /w:[ 9 ] /type:1
  //: joint g31 (CLR) @(485, 249) /w:[ -1 13 14 16 ]
  //: joint g22 (C) @(318, 137) /w:[ 20 22 -1 19 ]
  //: joint g98 (w6) @(528, 206) /w:[ 1 2 4 -1 ]
  //: LED g67 (w63) @(357,276) /sn:0 /w:[ 9 ] /type:1
  _GGAND2 #(6) g180 (.I0(w116), .I1(CLK), .Z(w40));   //: @(158,660) /sn:0 /w:[ 1 29 0 ]
  //: joint g99 (w63) @(523, 309) /w:[ 4 6 3 -1 ]
  //: joint g41 (w4) @(498, 259) /w:[ -1 10 20 9 ]
  //: joint g36 (w4) @(498, 665) /w:[ -1 2 28 1 ]
  //: joint g33 (CLR) @(485, 446) /w:[ -1 21 22 24 ]
  //: IN g45 (Add_A) @(567,-360) /sn:0 /R:3 /w:[ 0 ]
  //: IN g54 (rc_s) @(8,-204) /sn:0 /w:[ 0 ]
  //: joint g42 (w4) @(498, 164) /w:[ -1 12 18 11 ]
  //: LED g69 (w21) @(357,467) /sn:0 /w:[ 9 ] /type:1
  //: joint g40 (w4) @(498, 359) /w:[ -1 8 22 7 ]
  //: IN g52 (Add_B) @(673,-317) /sn:0 /R:3 /w:[ 0 ]
  _GGDECODER8 #(6, 6) g167 (.I(Add_A), .E(ra_s), .Z0(w27), .Z1(w31), .Z2(w34), .Z3(w39), .Z4(w46), .Z5(w53), .Z6(w59), .Z7(w65));   //: @(567,-258) /sn:0 /w:[ 1 1 1 1 0 0 0 0 0 0 ] /ss:0 /do:0
  //: LED g66 (w6) @(357,177) /sn:0 /w:[ 9 ] /type:1
  _GGBUFIF8 #(4, 6) g12 (.Z(B), .I(w23), .E(w55));   //: @(535,-8) /sn:0 /w:[ 9 5 1 ]
  //: joint g108 (A) @(705, 453) /w:[ -1 21 22 24 ]
  //: joint g46 (B) @(650, 309) /w:[ -1 4 14 3 ]
  //: joint g34 (CLR) @(485, 552) /w:[ -1 25 26 28 ]
  //: joint g28 (CLR) @(485, -58) /w:[ -1 2 1 4 ]
  //: joint g106 (A) @(705, 263) /w:[ -1 4 14 3 ]
  _GGBUFIF8 #(4, 6) g14 (.Z(B), .I(w6), .E(w61));   //: @(546,206) /sn:0 /w:[ 13 0 1 ]
  _GGREG8 #(10, 10, 20) g5 (.Q(w21), .D(C), .EN(w4), .CLR(~CLR), .CK(w25));   //: @(427,451) /sn:0 /w:[ 0 9 25 23 1 ]
  _GGAND2 #(6) g177 (.I0(w91), .I1(CLK), .Z(w20));   //: @(158,354) /sn:0 /w:[ 1 19 0 ]
  //: OUT g11 (B) @(862,379) /sn:0 /w:[ 0 ]
  //: joint g96 (w23) @(524, -8) /w:[ 4 6 3 -1 ]
  //: joint g187 (CLK) @(134, 453) /w:[ 22 21 -1 24 ]
  _GGBUFIF8 #(4, 6) g19 (.Z(B), .I(w36), .E(w76));   //: @(552,725) /sn:0 /w:[ 29 5 1 ]
  //: IN g21 (Add_C) @(96,-337) /sn:0 /R:3 /w:[ 0 ]
  //: joint g20 (C) @(318, 24) /w:[ 24 26 -1 23 ]
  //: joint g32 (CLR) @(485, 349) /w:[ -1 17 18 20 ]
  //: joint g78 (w72) @(429, 602) /w:[ 2 1 8 -1 ]
  //: joint g97 (w1) @(528, 92) /w:[ 1 2 4 -1 ]
  _GGAND2 #(6) g175 (.I0(w101), .I1(CLK), .Z(w10));   //: @(158,159) /sn:0 /w:[ 1 11 0 ]
  _GGAND2 #(6) g176 (.I0(w104), .I1(CLK), .Z(w15));   //: @(158,254) /sn:0 /w:[ 1 15 0 ]
  _GGBUFIF8 #(4, 6) g93 (.Z(A), .I(w21), .E(w53));   //: @(546,453) /sn:0 /w:[ 23 7 1 ]
  //: joint g100 (w16) @(519, 400) /w:[ 4 6 3 -1 ]
  //: joint g105 (A) @(705, 159) /w:[ -1 6 12 5 ]
  _GGBUFIF8 #(4, 6) g15 (.Z(B), .I(w63), .E(w64));   //: @(546,309) /sn:0 /w:[ 15 5 1 ]
  _GGBUFIF8 #(4, 6) g89 (.Z(A), .I(w1), .E(w31));   //: @(546,45) /sn:0 /w:[ 11 3 0 ]
  //: joint g38 (w4) @(498, 562) /w:[ -1 4 26 3 ]
  //: joint g43 (w4) @(498, 54) /w:[ -1 14 16 13 ]
  //: joint g101 (w21) @(522, 493) /w:[ 4 6 3 -1 ]
  //: joint g0 (A) @(705, 279) /w:[ 1 2 -1 16 ]
  //: joint g27 (C) @(318, 645) /w:[ 1 2 -1 28 ]
  //: joint g48 (B) @(650, 493) /w:[ -1 21 22 24 ]
  //: joint g171 (w23) @(421, -8) /w:[ 2 1 8 -1 ]
  //: joint g37 (B) @(650, 92) /w:[ -1 8 10 7 ]
  _GGBUFIF8 #(4, 6) g88 (.Z(A), .I(w23), .E(w27));   //: @(525,-59) /sn:0 /w:[ 9 7 0 ]
  _GGBUFIF8 #(4, 6) g95 (.Z(A), .I(w36), .E(w65));   //: @(552,685) /sn:0 /w:[ 29 7 1 ]
  //: IN g55 (CLR) @(460,-217) /sn:0 /R:2 /w:[ 3 ]
  _GGBUFIF8 #(4, 6) g13 (.Z(B), .I(w1), .E(w58));   //: @(546,92) /sn:0 /w:[ 11 0 1 ]
  //: joint g76 (w16) @(427, 400) /w:[ 2 1 8 -1 ]
  //: IN g53 (rb_s) @(602,-330) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin comparator
module comparator();
//: interface  /sz:(216, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls


endmodule
//: /netlistEnd

//: /netlistBegin sub_8
module sub_8(A, s, cout, B);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:1138,138)(1119,138)(1119,138)(1100,138){1}
//: {2}(1099,138)(968,138){3}
//: {4}(967,138)(831,138){5}
//: {6}(830,138)(698,138){7}
//: {8}(697,138)(560,138){9}
//: {10}(559,138)(490,138)(490,138)(421,138){11}
//: {12}(420,138)(287,138){13}
//: {14}(286,138)(143,138){15}
//: {16}(142,138)(3,138){17}
reg w7;    //: /sn:0 {0}(292,258)(292,180){1}
//: {2}(294,178)(424,178){3}
//: {4}(428,178)(496,178)(496,178)(563,178){5}
//: {6}(567,178)(635,178)(635,178)(702,178){7}
//: {8}(706,178)(770,178)(770,178)(834,178){9}
//: {10}(838,178)(905,178)(905,178)(971,178){11}
//: {12}(975,178)(1103,178){13}
//: {14}(1107,178)(1194,178){15}
//: {16}(1198,178)(1249,178){17}
//: {18}(1196,180)(1196,190)(1197,190)(1197,271){19}
//: {20}(1105,180)(1105,258){21}
//: {22}(973,180)(973,258){23}
//: {24}(836,180)(836,190)(836,190)(836,258){25}
//: {26}(704,180)(704,190)(704,190)(704,258){27}
//: {28}(565,180)(565,190)(565,190)(565,258){29}
//: {30}(426,180)(426,258){31}
//: {32}(290,178)(150,178){33}
//: {34}(146,178)(13,178)(13,365)(17,365){35}
//: {36}(19,363)(19,356){37}
//: {38}(19,367)(19,375){39}
//: {40}(148,180)(148,219)(149,219)(149,258){41}
input [7:0] A;    //: /sn:0 {0}(#:1138,99)(1063,99){1}
//: {2}(1062,99)(933,99){3}
//: {4}(932,99)(795,99){5}
//: {6}(794,99)(658,99){7}
//: {8}(657,99)(521,99){9}
//: {10}(520,99)(382,99){11}
//: {12}(381,99)(251,99){13}
//: {14}(250,99)(106,99){15}
//: {16}(105,99)(4,99){17}
reg w12;    //: /sn:0 {0}(1153,237)(1153,241)(1192,241)(1192,271){1}
output [7:0] s;    //: /sn:0 {0}(620,393)(#:620,460){1}
output cout;    //: /sn:0 {0}(21,396)(21,410)(38,410){1}
wire w16;    //: /sn:0 {0}(658,103)(658,111)(661,111)(661,324){1}
wire w13;    //: /sn:0 {0}(775,356)(735,356){1}
wire w6;    //: /sn:0 {0}(933,103)(933,111)(931,111)(931,328){1}
wire w50;    //: /sn:0 {0}(421,142)(421,258){1}
wire w34;    //: /sn:0 {0}(275,384)(275,484)(595,484)(595,466){1}
wire w4;    //: /sn:0 {0}(655,466)(655,476)(1090,476)(1090,396){1}
wire w25;    //: /sn:0 {0}(423,320)(423,279){1}
wire w39;    //: /sn:0 {0}(132,382)(132,478)(585,478)(585,466){1}
wire w56;    //: /sn:0 {0}(143,142)(143,200)(144,200)(144,258){1}
wire w22;    //: /sn:0 {0}(549,388)(549,497)(615,497)(615,466){1}
wire w36;    //: /sn:0 {0}(106,103)(106,316){1}
wire w0;    //: /sn:0 {0}(1102,279)(1102,315)(1104,315)(1104,330){1}
wire w3;    //: /sn:0 {0}(1043,360)(1023,360)(1023,360)(1005,360){1}
wire w20;    //: /sn:0 {0}(562,279)(562,307)(563,307)(563,322){1}
wire w30;    //: /sn:0 {0}(289,279)(289,318){1}
wire w29;    //: /sn:0 {0}(409,386)(409,491)(605,491)(605,466){1}
wire w18;    //: /sn:0 {0}(640,354)(612,354)(612,354)(597,354){1}
wire w19;    //: /sn:0 {0}(687,390)(687,496)(625,496)(625,466){1}
wire w23;    //: /sn:0 {0}(502,352)(457,352){1}
wire w10;    //: /sn:0 {0}(833,279)(833,302)(836,302)(836,326){1}
wire w21;    //: /sn:0 {0}(521,103)(521,111)(523,111)(523,322){1}
wire w31;    //: /sn:0 {0}(251,103)(251,111)(249,111)(249,318){1}
wire w1;    //: /sn:0 {0}(1063,103)(1063,111)(1064,111)(1064,330){1}
wire w32;    //: /sn:0 {0}(968,142)(968,258){1}
wire w53;    //: /sn:0 {0}(287,142)(287,258){1}
wire w8;    //: /sn:0 {0}(910,358)(870,358){1}
wire w44;    //: /sn:0 {0}(698,142)(698,200)(699,200)(699,258){1}
wire w17;    //: /sn:0 {0}(1100,142)(1100,150)(1100,150)(1100,258){1}
wire w35;    //: /sn:0 {0}(146,279)(146,308)(146,308)(146,316){1}
wire w28;    //: /sn:0 {0}(362,350)(323,350){1}
wire w33;    //: /sn:0 {0}(228,348)(195,348)(195,348)(180,348){1}
wire w14;    //: /sn:0 {0}(822,392)(822,488)(635,488)(635,466){1}
wire w11;    //: /sn:0 {0}(795,103)(795,111)(796,111)(796,326){1}
wire w2;    //: /sn:0 {0}(1194,292)(1194,362)(1138,362){1}
wire w41;    //: /sn:0 {0}(831,142)(831,258){1}
wire w47;    //: /sn:0 {0}(560,142)(560,200)(560,200)(560,258){1}
wire w15;    //: /sn:0 {0}(701,279)(701,324){1}
wire w38;    //: /sn:0 {0}(85,346)(24,346)(24,375){1}
wire w5;    //: /sn:0 {0}(970,279)(970,313)(971,313)(971,328){1}
wire w26;    //: /sn:0 {0}(382,103)(382,111)(383,111)(383,320){1}
wire w9;    //: /sn:0 {0}(957,394)(957,481)(645,481)(645,466){1}
//: enddecls

  F_Add g4 (.a(w21), .b(w20), .cin(w18), .cout(w23), .sum(w22));   //: @(503, 323) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: IN g8 (A) @(1140,99) /sn:0 /R:2 /w:[ 0 ]
  assign w56 = B[7]; //: TAP g44 @(143,136) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  F_Add g3 (.a(w16), .b(w15), .cin(w13), .cout(w18), .sum(w19));   //: @(641, 325) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w36 = A[7]; //: TAP g16 @(106,97) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  //: DIP g47 (w12) @(1153,227) /sn:0 /w:[ 0 ] /st:0 /dn:1
  assign w31 = A[6]; //: TAP g17 @(251,97) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  _GGXOR2 #(8) g26 (.I0(w7), .I1(w56), .Z(w35));   //: @(146,269) /sn:0 /R:3 /w:[ 41 1 0 ]
  F_Add g2 (.a(w11), .b(w10), .cin(w8), .cout(w13), .sum(w14));   //: @(776, 327) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  _GGXOR2 #(8) g23 (.I0(w7), .I1(w47), .Z(w20));   //: @(562,269) /sn:0 /R:3 /w:[ 29 1 0 ]
  //: joint g30 (w7) @(292, 178) /w:[ 2 -1 32 1 ]
  F_Add g1 (.a(w1), .b(w0), .cin(w2), .cout(w3), .sum(w4));   //: @(1044, 331) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  _GGXOR2 #(8) g24 (.I0(w7), .I1(w50), .Z(w25));   //: @(423,269) /sn:0 /R:3 /w:[ 31 1 1 ]
  assign w41 = B[2]; //: TAP g39 @(831,136) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: joint g29 (w7) @(148, 178) /w:[ 33 -1 34 40 ]
  //: SWITCH g18 (w7) @(1267,178) /sn:0 /R:2 /w:[ 17 ] /st:1 /dn:1
  assign w1 = A[0]; //: TAP g10 @(1063,97) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  _GGXOR2 #(8) g25 (.I0(w7), .I1(w53), .Z(w30));   //: @(289,269) /sn:0 /R:3 /w:[ 0 1 0 ]
  //: OUT g49 (s) @(620,396) /sn:0 /R:1 /w:[ 0 ]
  F_Add g6 (.a(w31), .b(w30), .cin(w28), .cout(w33), .sum(w34));   //: @(229, 319) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: OUT g50 (cout) @(35,410) /sn:0 /w:[ 1 ]
  F_Add g7 (.a(w36), .b(w35), .cin(w33), .cout(w38), .sum(w39));   //: @(86, 317) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: IN g9 (B) @(1140,138) /sn:0 /R:2 /w:[ 0 ]
  //: joint g35 (w7) @(973, 178) /w:[ 12 -1 11 22 ]
  _GGXOR2 #(8) g22 (.I0(w7), .I1(w44), .Z(w15));   //: @(701,269) /sn:0 /R:3 /w:[ 27 1 0 ]
  //: joint g31 (w7) @(565, 178) /w:[ 6 -1 5 28 ]
  //: joint g33 (w7) @(704, 178) /w:[ 8 -1 7 26 ]
  //: joint g36 (w7) @(836, 178) /w:[ 10 -1 9 24 ]
  assign w47 = B[4]; //: TAP g41 @(560,136) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  //: joint g45 (w7) @(19, 365) /w:[ -1 36 35 38 ]
  assign w44 = B[3]; //: TAP g40 @(698,136) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  assign w50 = B[5]; //: TAP g42 @(421,136) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  assign w11 = A[2]; //: TAP g12 @(795,97) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  _GGXOR2 #(8) g28 (.I0(w38), .I1(w7), .Z(cout));   //: @(21,386) /sn:0 /R:3 /w:[ 1 39 0 ]
  //: joint g34 (w7) @(1105, 178) /w:[ 14 -1 13 20 ]
  //: joint g46 (w7) @(1196, 178) /w:[ 16 -1 15 18 ]
  F_Add g5 (.a(w26), .b(w25), .cin(w23), .cout(w28), .sum(w29));   //: @(363, 321) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  assign w6 = A[1]; //: TAP g11 @(933,97) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  assign w21 = A[4]; //: TAP g14 @(521,97) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  _GGXOR2 #(8) g19 (.I0(w7), .I1(w17), .Z(w0));   //: @(1102,269) /sn:0 /R:3 /w:[ 21 1 0 ]
  _GGXOR2 #(8) g21 (.I0(w7), .I1(w41), .Z(w10));   //: @(833,269) /sn:0 /R:3 /w:[ 25 1 0 ]
  _GGXOR2 #(8) g20 (.I0(w7), .I1(w32), .Z(w5));   //: @(970,269) /sn:0 /R:3 /w:[ 23 1 0 ]
  //: joint g32 (w7) @(426, 178) /w:[ 4 -1 3 30 ]
  F_Add g0 (.a(w6), .b(w5), .cin(w3), .cout(w8), .sum(w9));   //: @(911, 329) /sz:(93, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w26 = A[5]; //: TAP g15 @(382,97) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  assign w32 = B[1]; //: TAP g38 @(968,136) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  assign w53 = B[6]; //: TAP g43 @(287,136) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  _GGXOR2 #(8) g27 (.I0(w7), .I1(w12), .Z(w2));   //: @(1194,282) /sn:0 /R:3 /w:[ 19 1 0 ]
  assign s = {w39, w34, w29, w22, w19, w14, w9, w4}; //: CONCAT g48  @(620,461) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 0 ] /dr:0 /tp:0 /drp:1
  assign w17 = B[0]; //: TAP g37 @(1100,136) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  assign w16 = A[3]; //: TAP g13 @(658,97) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1

endmodule
//: /netlistEnd

